<?xml version="1.0" encoding="ISO-8859-1"?>
<!DOCTYPE svg PUBLIC '-//W3C//DTD SVG 1.0//EN'
          'http://www.w3.org/TR/2001/REC-SVG-20010904/DTD/svg10.dtd'>
<svg xmlns:xlink="http://www.w3.org/1999/xlink" style="fill-opacity:1; color-rendering:auto; color-interpolation:auto; text-rendering:auto; stroke:black; stroke-linecap:square; stroke-miterlimit:10; shape-rendering:auto; stroke-opacity:1; fill:black; stroke-dasharray:none; font-weight:normal; stroke-width:1; font-family:'Dialog'; font-style:normal; stroke-linejoin:miter; font-size:12px; stroke-dashoffset:0; image-rendering:auto;" width="1920" height="1080" xmlns="http://www.w3.org/2000/svg"
><!--Generated by the Batik Graphics2D SVG Generator--><defs id="genericDefs"
  /><g
  ><g style="stroke-width:0.2;"
    ><path style="fill:none;" d="M479.43 132.99 L439.04 147.17 L430.66 165.82 L431.39 167.69 L470.27 187.93 L499.24 166.04 L499.05 151.69 L479.43 132.99 Z"
      /><path d="M479.43 132.99 L439.04 147.17 L430.66 165.82 L431.39 167.69 L470.27 187.93 L499.24 166.04 L499.05 151.69 L479.43 132.99 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M949.71 24.77 L922.97 38.36 L919.69 53.37 L933.02 72.36 L969.87 62.79 L975.05 56.27 L949.71 24.77 Z"
      /><path d="M949.71 24.77 L922.97 38.36 L919.69 53.37 L933.02 72.36 L969.87 62.79 L975.05 56.27 L949.71 24.77 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1563.17 322.56 L1585.96 348.11 L1576.59 378.5 L1541.99 380.52 L1524.1899 355.32 L1531.12 332.34 L1563.17 322.56 Z"
      /><path d="M1563.17 322.56 L1585.96 348.11 L1576.59 378.5 L1541.99 380.52 L1524.1899 355.32 L1531.12 332.34 L1563.17 322.56 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1694.37 815.1 L1682.53 844.74 L1648.99 842.56 L1639.54 813.74 L1664.6899 792.94 L1694.37 815.1 Z"
      /><path d="M1694.37 815.1 L1682.53 844.74 L1648.99 842.56 L1639.54 813.74 L1664.6899 792.94 L1694.37 815.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M149.63 603.43 L177.28 610.31 L173.21 653.57 L146.23 666.74 L143.06 665.78 L124.92 627.38 L149.63 603.43 Z"
      /><path d="M149.63 603.43 L177.28 610.31 L173.21 653.57 L146.23 666.74 L143.06 665.78 L124.92 627.38 L149.63 603.43 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1684.7 0 L1695.16 51.68 L1684.61 63.43 L1646.73 59.3 L1640.55 49.3 L1653 0 L1684.7 0 Z"
      /><path d="M1684.7 0 L1695.16 51.68 L1684.61 63.43 L1646.73 59.3 L1640.55 49.3 L1653 0 L1684.7 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1637.89 423.52 L1616.85 443.42 L1624.72 481.14 L1667.64 468.75 L1671.58 435.08 L1637.89 423.52 Z"
      /><path d="M1637.89 423.52 L1616.85 443.42 L1624.72 481.14 L1667.64 468.75 L1671.58 435.08 L1637.89 423.52 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M813.29 253.07 L805.24 244.96 L762.93 247.53 L752.48 261.1 L752.9 269.91 L790.1 300.51 L806.07 297.96 L813.29 253.07 Z"
      /><path d="M813.29 253.07 L805.24 244.96 L762.93 247.53 L752.48 261.1 L752.9 269.91 L790.1 300.51 L806.07 297.96 L813.29 253.07 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1340.75 119.08 L1317.6899 119.5 L1298.36 142.34 L1312.6 172.23 L1343.85 166.16 L1349.73 128.01 L1340.75 119.08 Z"
      /><path d="M1340.75 119.08 L1317.6899 119.5 L1298.36 142.34 L1312.6 172.23 L1343.85 166.16 L1349.73 128.01 L1340.75 119.08 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1549.3101 924.65 L1527.22 935.08 L1522.3 971.41 L1552.85 991.24 L1580.3 948.58 L1576.95 937.25 L1549.3101 924.65 Z"
      /><path d="M1549.3101 924.65 L1527.22 935.08 L1522.3 971.41 L1552.85 991.24 L1580.3 948.58 L1576.95 937.25 L1549.3101 924.65 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1407.6899 435.48 L1365.66 422.98 L1359.45 428.61 L1353.6801 457.3 L1386.13 484.95 L1409.78 472.26 L1407.6899 435.48 Z"
      /><path d="M1407.6899 435.48 L1365.66 422.98 L1359.45 428.61 L1353.6801 457.3 L1386.13 484.95 L1409.78 472.26 L1407.6899 435.48 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M728.43 904.21 L710.43 928.48 L727.4 954.25 L766.93 949.45 L773 939.25 L761.68 907.08 L728.43 904.21 Z"
      /><path d="M728.43 904.21 L710.43 928.48 L727.4 954.25 L766.93 949.45 L773 939.25 L761.68 907.08 L728.43 904.21 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M962.25 174.19 L990.28 191.51 L985.61 219.15 L939.82 209.71 L962.25 174.19 Z"
      /><path d="M962.25 174.19 L990.28 191.51 L985.61 219.15 L939.82 209.71 L962.25 174.19 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1814.54 756.59 L1804.4301 763.91 L1801.16 803.13 L1830.84 815.43 L1857.22 787.4 L1839.4 759.4 L1814.54 756.59 Z"
      /><path d="M1814.54 756.59 L1804.4301 763.91 L1801.16 803.13 L1830.84 815.43 L1857.22 787.4 L1839.4 759.4 L1814.54 756.59 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1758.04 536.89 L1721.35 529.12 L1706.4301 541.91 L1712.83 573.46 L1743.5699 581.99 L1748.92 579.08 L1760.2 541.89 L1758.04 536.89 Z"
      /><path d="M1758.04 536.89 L1721.35 529.12 L1706.4301 541.91 L1712.83 573.46 L1743.5699 581.99 L1748.92 579.08 L1760.2 541.89 L1758.04 536.89 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M376.77 1045.8199 L339.26 1030.47 L319.62 1049.8199 L320.2 1080 L377.8 1080 L376.77 1045.8199 Z"
      /><path d="M376.77 1045.8199 L339.26 1030.47 L319.62 1049.8199 L320.2 1080 L377.8 1080 L376.77 1045.8199 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M209.56 30.24 L177.13 47.26 L184.03 81.23 L198.32 86.07 L231.27 63.19 L231.98 51.27 L209.56 30.24 Z"
      /><path d="M209.56 30.24 L177.13 47.26 L184.03 81.23 L198.32 86.07 L231.27 63.19 L231.98 51.27 L209.56 30.24 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M282.77 431.58 L259.37 411.88 L236.9 414.18 L223.86 448.02 L232.17 464.38 L268.31 469.82 L282.39 453.74 L282.77 431.58 Z"
      /><path d="M282.77 431.58 L259.37 411.88 L236.9 414.18 L223.86 448.02 L232.17 464.38 L268.31 469.82 L282.39 453.74 L282.77 431.58 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M772.5 795.16 L812.16 818.03 L807.25 836.89 L768.11 851.21 L754.18 816.75 L772.5 795.16 Z"
      /><path d="M772.5 795.16 L812.16 818.03 L807.25 836.89 L768.11 851.21 L754.18 816.75 L772.5 795.16 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M955.65 935.97 L921.95 936.04 L914.2 944.68 L915.26 970.5 L941.18 993.83 L973.36 970.28 L955.65 935.97 Z"
      /><path d="M955.65 935.97 L921.95 936.04 L914.2 944.68 L915.26 970.5 L941.18 993.83 L973.36 970.28 L955.65 935.97 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1173.71 558.86 L1213.5 583.27 L1191.1899 614.86 L1166.3 613.19 L1151.22 582 L1173.71 558.86 Z"
      /><path d="M1173.71 558.86 L1213.5 583.27 L1191.1899 614.86 L1166.3 613.19 L1151.22 582 L1173.71 558.86 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M397.76 839.54 L367.78 832.42 L345.55 869.3 L367.83 885.59 L397.9 871.63 L397.76 839.54 Z"
      /><path d="M397.76 839.54 L367.78 832.42 L345.55 869.3 L367.83 885.59 L397.9 871.63 L397.76 839.54 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M288.56 228.92 L259.4 235.26 L251.51 257.39 L278.6 277.5 L287.48 275.3 L302.9 240.59 L288.56 228.92 Z"
      /><path d="M288.56 228.92 L259.4 235.26 L251.51 257.39 L278.6 277.5 L287.48 275.3 L302.9 240.59 L288.56 228.92 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M851.3 0 L851.97 34.74 L815.66 40.29 L812.4 36.93 L815 0 L851.3 0 Z"
      /><path d="M851.3 0 L851.97 34.74 L815.66 40.29 L812.4 36.93 L815 0 L851.3 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1125.02 634.37 L1147.48 636.09 L1164.4399 669.08 L1144.88 689.96 L1104.9399 675.44 L1102.67 667.12 L1125.02 634.37 Z"
      /><path d="M1125.02 634.37 L1147.48 636.09 L1164.4399 669.08 L1144.88 689.96 L1104.9399 675.44 L1102.67 667.12 L1125.02 634.37 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1809.04 711.71 L1814.54 756.59 L1804.4301 763.91 L1765.52 753.44 L1763.97 730.85 L1792.45 707.66 L1809.04 711.71 Z"
      /><path d="M1809.04 711.71 L1814.54 756.59 L1804.4301 763.91 L1765.52 753.44 L1763.97 730.85 L1792.45 707.66 L1809.04 711.71 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M948.88 824.39 L980.08 830.88 L989 857.11 L954.76 881.86 L945.38 879.16 L931.61 843.01 L948.88 824.39 Z"
      /><path d="M948.88 824.39 L980.08 830.88 L989 857.11 L954.76 881.86 L945.38 879.16 L931.61 843.01 L948.88 824.39 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M334.9 151.1 L305.2 114.94 L275.98 132.95 L279.8 154.9 L317.62 169.04 L334.9 151.1 Z"
      /><path d="M334.9 151.1 L305.2 114.94 L275.98 132.95 L279.8 154.9 L317.62 169.04 L334.9 151.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M947.36 369.3 L920.81 399.33 L899.98 393.03 L895.63 356.02 L929.17 343.39 L947.36 369.3 Z"
      /><path d="M947.36 369.3 L920.81 399.33 L899.98 393.03 L895.63 356.02 L929.17 343.39 L947.36 369.3 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M98.03 150.45 L110.36 177.97 L92.46 196.84 L72.29 195.66 L63.76 161.34 L98.03 150.45 Z"
      /><path d="M98.03 150.45 L110.36 177.97 L92.46 196.84 L72.29 195.66 L63.76 161.34 L98.03 150.45 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M603.85 93.07 L589.47 105.36 L589.86 140.28 L621.14 154.44 L638.35 145.03 L642.32 100.73 L634.78 93.96 L603.85 93.07 Z"
      /><path d="M603.85 93.07 L589.47 105.36 L589.86 140.28 L621.14 154.44 L638.35 145.03 L642.32 100.73 L634.78 93.96 L603.85 93.07 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M897.5 0 L898.41 12.65 L922.97 38.36 L949.71 24.77 L954.6 0 L897.5 0 Z"
      /><path d="M897.5 0 L898.41 12.65 L922.97 38.36 L949.71 24.77 L954.6 0 L897.5 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1682.29 236.85 L1697.9 243.59 L1705.99 265.71 L1692.26 288.19 L1665.37 291.54 L1650.98 275.8 L1654.2 246.08 L1682.29 236.85 Z"
      /><path d="M1682.29 236.85 L1697.9 243.59 L1705.99 265.71 L1692.26 288.19 L1665.37 291.54 L1650.98 275.8 L1654.2 246.08 L1682.29 236.85 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M765.86 451.7 L759.85 474.33 L734.69 487.02 L712.24 461.71 L719.69 431.88 L737.98 427.65 L765.86 451.7 Z"
      /><path d="M765.86 451.7 L759.85 474.33 L734.69 487.02 L712.24 461.71 L719.69 431.88 L737.98 427.65 L765.86 451.7 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1712.83 573.46 L1694.01 590.7 L1694.23 600.99 L1715.5699 622.87 L1736.39 621.14 L1743.5699 581.99 L1712.83 573.46 Z"
      /><path d="M1712.83 573.46 L1694.01 590.7 L1694.23 600.99 L1715.5699 622.87 L1736.39 621.14 L1743.5699 581.99 L1712.83 573.46 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M947.36 369.3 L968.88 372.04 L975.92 380.31 L969.66 418.72 L933.12 420.38 L920.81 399.33 L947.36 369.3 Z"
      /><path d="M947.36 369.3 L968.88 372.04 L975.92 380.31 L969.66 418.72 L933.12 420.38 L920.81 399.33 L947.36 369.3 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1009.14 429.87 L1024 447.36 L1005.05 483.78 L966.19 472.72 L979.53 429.52 L1009.14 429.87 Z"
      /><path d="M1009.14 429.87 L1024 447.36 L1005.05 483.78 L966.19 472.72 L979.53 429.52 L1009.14 429.87 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M1530.03 879.33 L1548.49 890.21 L1549.3101 924.65 L1527.22 935.08 L1500.26 919.25 L1503.55 889.62 L1530.03 879.33 Z"
      /><path d="M1530.03 879.33 L1548.49 890.21 L1549.3101 924.65 L1527.22 935.08 L1500.26 919.25 L1503.55 889.62 L1530.03 879.33 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M397.99 245.7 L372.4 256.04 L372.4 278.7 L395.27 299.37 L418.45 287.56 L421.8 265.31 L397.99 245.7 Z"
      /><path d="M397.99 245.7 L372.4 256.04 L372.4 278.7 L395.27 299.37 L418.45 287.56 L421.8 265.31 L397.99 245.7 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M848.78 250.57 L813.29 253.07 L806.07 297.96 L820.14 307.27 L843.69 303.41 L861.05 276.9 L848.78 250.57 Z"
      /><path d="M848.78 250.57 L813.29 253.07 L806.07 297.96 L820.14 307.27 L843.69 303.41 L861.05 276.9 L848.78 250.57 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M553.34 428.25 L571.04 434.9 L581.12 475.22 L558.18 491.95 L545.94 491.11 L530.85 475.57 L536.26 437.55 L553.34 428.25 Z"
      /><path d="M553.34 428.25 L571.04 434.9 L581.12 475.22 L558.18 491.95 L545.94 491.11 L530.85 475.57 L536.26 437.55 L553.34 428.25 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M523.99 523.57 L546.29 553.73 L523.98 572.82 L491.54 564.82 L486.4 551.71 L501.97 523.26 L523.99 523.57 Z"
      /><path d="M523.99 523.57 L546.29 553.73 L523.98 572.82 L491.54 564.82 L486.4 551.71 L501.97 523.26 L523.99 523.57 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M540.59 663.3 L563.86 696.82 L543.72 724.37 L524.87 719.02 L510.79 685.97 L523.19 667.27 L540.59 663.3 Z"
      /><path d="M540.59 663.3 L563.86 696.82 L543.72 724.37 L524.87 719.02 L510.79 685.97 L523.19 667.27 L540.59 663.3 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1028.23 645.64 L1050.76 657.78 L1047.13 701.58 L996.81 691 L991.48 681.3 L993.99 670.18 L1028.23 645.64 Z"
      /><path d="M1028.23 645.64 L1050.76 657.78 L1047.13 701.58 L996.81 691 L991.48 681.3 L993.99 670.18 L1028.23 645.64 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M411.99 829.27 L397.76 839.54 L397.9 871.63 L418.35 886.73 L443.67 875.98 L448.19 851.13 L411.99 829.27 Z"
      /><path d="M411.99 829.27 L397.76 839.54 L397.9 871.63 L418.35 886.73 L443.67 875.98 L448.19 851.13 L411.99 829.27 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M910.74 750.48 L885.39 735.96 L859.86 756.17 L872.13 789.82 L900.09 794.63 L907.04 789.93 L910.74 750.48 Z"
      /><path d="M910.74 750.48 L885.39 735.96 L859.86 756.17 L872.13 789.82 L900.09 794.63 L907.04 789.93 L910.74 750.48 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1270.09 97.69 L1254.01 95.75 L1232.78 128.19 L1258.83 150.29 L1279 138.59 L1270.09 97.69 Z"
      /><path d="M1270.09 97.69 L1254.01 95.75 L1232.78 128.19 L1258.83 150.29 L1279 138.59 L1270.09 97.69 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M996.58 282.81 L1014.29 297.03 L1008.16 332.35 L982.07 334.86 L966.56 319.17 L970.15 296.5 L996.58 282.81 Z"
      /><path d="M996.58 282.81 L1014.29 297.03 L1008.16 332.35 L982.07 334.86 L966.56 319.17 L970.15 296.5 L996.58 282.81 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M35.38 359.87 L0 363.9 L0 410.6 L43.42 401.24 L47.09 371.1 L35.38 359.87 Z"
      /><path d="M35.38 359.87 L0 363.9 L0 410.6 L43.42 401.24 L47.09 371.1 L35.38 359.87 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1013.26 177.72 L1034.9301 207.71 L1022.59 227.53 L985.66 219.24 L985.61 219.15 L990.28 191.51 L1013.26 177.72 Z"
      /><path d="M1013.26 177.72 L1034.9301 207.71 L1022.59 227.53 L985.66 219.24 L985.61 219.15 L990.28 191.51 L1013.26 177.72 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M107.18 683.97 L79.12 653.1 L56.62 654.41 L51.3 659.49 L51.3 709.24 L91.58 717.52 L101.48 710.87 L107.18 683.97 Z"
      /><path d="M107.18 683.97 L79.12 653.1 L56.62 654.41 L51.3 659.49 L51.3 709.24 L91.58 717.52 L101.48 710.87 L107.18 683.97 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1119.85 1053.75 L1107.83 1041.97 L1072.4 1052.15 L1069.2 1080 L1120.4 1080 L1119.85 1053.75 Z"
      /><path d="M1119.85 1053.75 L1107.83 1041.97 L1072.4 1052.15 L1069.2 1080 L1120.4 1080 L1119.85 1053.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1566.74 168.99 L1569.9 171.75 L1575.04 211.24 L1567.4399 219.02 L1537.74 219.4 L1531 214.44 L1529.48 194.77 L1550.15 170.6 L1566.74 168.99 Z"
      /><path d="M1566.74 168.99 L1569.9 171.75 L1575.04 211.24 L1567.4399 219.02 L1537.74 219.4 L1531 214.44 L1529.48 194.77 L1550.15 170.6 L1566.74 168.99 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M159.05 96.42 L158.14 99.31 L125.95 116.48 L102.67 88.94 L132.33 67.23 L159.05 96.42 Z"
      /><path d="M159.05 96.42 L158.14 99.31 L125.95 116.48 L102.67 88.94 L132.33 67.23 L159.05 96.42 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M36.19 290.19 L16.16 314.53 L38.53 333.85 L65.86 319.78 L64.57 301.08 L36.19 290.19 Z"
      /><path d="M36.19 290.19 L16.16 314.53 L38.53 333.85 L65.86 319.78 L64.57 301.08 L36.19 290.19 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1014.8 87.25 L1041.99 101.03 L1044.47 128.92 L1038 136.43 L990.54 119.73 L989.56 116.82 L1014.8 87.25 Z"
      /><path d="M1014.8 87.25 L1041.99 101.03 L1044.47 128.92 L1038 136.43 L990.54 119.73 L989.56 116.82 L1014.8 87.25 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1462.55 464.68 L1433.5699 482.78 L1438.78 514.74 L1458.8101 525.16 L1491.87 506.53 L1492.12 488.01 L1462.55 464.68 Z"
      /><path d="M1462.55 464.68 L1433.5699 482.78 L1438.78 514.74 L1458.8101 525.16 L1491.87 506.53 L1492.12 488.01 L1462.55 464.68 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M990.54 119.73 L1038 136.43 L1035.97 154.78 L1014.77 171.79 L985.09 143.44 L990.54 119.73 Z"
      /><path d="M990.54 119.73 L1038 136.43 L1035.97 154.78 L1014.77 171.79 L985.09 143.44 L990.54 119.73 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1147.16 714.99 L1107.9301 734.61 L1105.23 743.89 L1126.45 772.08 L1162.52 763.16 L1168.15 731.16 L1147.16 714.99 Z"
      /><path d="M1147.16 714.99 L1107.9301 734.61 L1105.23 743.89 L1126.45 772.08 L1162.52 763.16 L1168.15 731.16 L1147.16 714.99 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M917.04 1020.82 L887.54 1012.41 L875.24 1040.15 L900.49 1062.0699 L921.31 1041.76 L917.04 1020.82 Z"
      /><path d="M917.04 1020.82 L887.54 1012.41 L875.24 1040.15 L900.49 1062.0699 L921.31 1041.76 L917.04 1020.82 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1505.8 0 L1551.5 0 L1550.34 39 L1531.3101 51.27 L1504.71 36.89 L1505.8 0 Z"
      /><path d="M1505.8 0 L1551.5 0 L1550.34 39 L1531.3101 51.27 L1504.71 36.89 L1505.8 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M832.16 705.26 L801.92 679.22 L773.1 694.79 L770.25 716.02 L787.64 733.54 L826.4 722.82 L832.16 705.26 Z"
      /><path d="M832.16 705.26 L801.92 679.22 L773.1 694.79 L770.25 716.02 L787.64 733.54 L826.4 722.82 L832.16 705.26 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1166.3 613.19 L1191.1899 614.86 L1205.76 641.62 L1185.37 670.21 L1164.4399 669.08 L1147.48 636.09 L1166.3 613.19 Z"
      /><path d="M1166.3 613.19 L1191.1899 614.86 L1205.76 641.62 L1185.37 670.21 L1164.4399 669.08 L1147.48 636.09 L1166.3 613.19 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M118.72 953.85 L117.22 954.11 L92.85 991.55 L115.71 1030.67 L150.41 1017.44 L156.38 1005.65 L118.72 953.85 Z"
      /><path d="M118.72 953.85 L117.22 954.11 L92.85 991.55 L115.71 1030.67 L150.41 1017.44 L156.38 1005.65 L118.72 953.85 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M313.79 239.76 L332.99 254.75 L326.64 291.37 L317.91 294.11 L287.48 275.3 L302.9 240.59 L313.79 239.76 Z"
      /><path d="M313.79 239.76 L332.99 254.75 L326.64 291.37 L317.91 294.11 L287.48 275.3 L302.9 240.59 L313.79 239.76 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1104.9399 675.44 L1144.88 689.96 L1147.16 714.99 L1107.9301 734.61 L1090.24 701.39 L1104.9399 675.44 Z"
      /><path d="M1104.9399 675.44 L1144.88 689.96 L1147.16 714.99 L1107.9301 734.61 L1090.24 701.39 L1104.9399 675.44 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M787.64 733.54 L770.25 716.02 L733.93 731.16 L740.71 762.95 L772.3 775.8 L785.78 764.01 L787.64 733.54 Z"
      /><path d="M787.64 733.54 L770.25 716.02 L733.93 731.16 L740.71 762.95 L772.3 775.8 L785.78 764.01 L787.64 733.54 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M154.2 216.22 L139 210.26 L109.45 229.29 L106.32 239.18 L107.2 241.41 L142.03 261.28 L162.79 246.69 L154.2 216.22 Z"
      /><path d="M154.2 216.22 L139 210.26 L109.45 229.29 L106.32 239.18 L107.2 241.41 L142.03 261.28 L162.79 246.69 L154.2 216.22 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M462.3 0 L505.4 0 L504.72 43.19 L473.44 48.47 L458.44 25.86 L462.3 0 Z"
      /><path d="M462.3 0 L505.4 0 L504.72 43.19 L473.44 48.47 L458.44 25.86 L462.3 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M772.3 775.8 L772.5 795.16 L754.18 816.75 L726.71 813.38 L714.19 786.36 L740.71 762.95 L772.3 775.8 Z"
      /><path d="M772.3 775.8 L772.5 795.16 L754.18 816.75 L726.71 813.38 L714.19 786.36 L740.71 762.95 L772.3 775.8 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M907.04 789.93 L941.32 796.47 L948.88 824.39 L931.61 843.01 L900.52 839.99 L900.09 794.63 L907.04 789.93 Z"
      /><path d="M907.04 789.93 L941.32 796.47 L948.88 824.39 L931.61 843.01 L900.52 839.99 L900.09 794.63 L907.04 789.93 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M197.79 565.9 L190.14 550.37 L142.31 558.6 L135.95 570.82 L149.63 603.43 L177.28 610.31 L179.7 609.15 L197.79 565.9 Z"
      /><path d="M197.79 565.9 L190.14 550.37 L142.31 558.6 L135.95 570.82 L149.63 603.43 L177.28 610.31 L179.7 609.15 L197.79 565.9 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1792.45 707.66 L1763.97 730.85 L1739.62 713.88 L1746.17 679.46 L1777.33 678.61 L1792.45 707.66 Z"
      /><path d="M1792.45 707.66 L1763.97 730.85 L1739.62 713.88 L1746.17 679.46 L1777.33 678.61 L1792.45 707.66 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M385.14 368.51 L360.13 389.86 L362.87 413.88 L378.52 423 L409.03 410.13 L411.72 389.83 L385.14 368.51 Z"
      /><path d="M385.14 368.51 L360.13 389.86 L362.87 413.88 L378.52 423 L409.03 410.13 L411.72 389.83 L385.14 368.51 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1731.4 0 L1684.7 0 L1695.16 51.68 L1730.49 49.14 L1737.02 40.24 L1731.4 0 Z"
      /><path d="M1731.4 0 L1684.7 0 L1695.16 51.68 L1730.49 49.14 L1737.02 40.24 L1731.4 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1759.11 159.24 L1754.21 172.13 L1710.73 178.37 L1704.8199 146.48 L1735.51 125.18 L1759.11 159.24 Z"
      /><path d="M1759.11 159.24 L1754.21 172.13 L1710.73 178.37 L1704.8199 146.48 L1735.51 125.18 L1759.11 159.24 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1667.64 468.75 L1685.23 487.01 L1668.86 521.26 L1641.65 517.77 L1623.87 482.73 L1624.72 481.14 L1667.64 468.75 Z"
      /><path d="M1667.64 468.75 L1685.23 487.01 L1668.86 521.26 L1641.65 517.77 L1623.87 482.73 L1624.72 481.14 L1667.64 468.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1232.78 128.19 L1258.83 150.29 L1253.75 172.39 L1221.03 181.57 L1205.48 143.66 L1216.8 129.24 L1232.78 128.19 Z"
      /><path d="M1232.78 128.19 L1258.83 150.29 L1253.75 172.39 L1221.03 181.57 L1205.48 143.66 L1216.8 129.24 L1232.78 128.19 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1139.72 294.11 L1118.59 263.76 L1089.85 272.08 L1082.46 298.65 L1101.7 317.62 L1136.0699 308.24 L1139.72 294.11 Z"
      /><path d="M1139.72 294.11 L1118.59 263.76 L1089.85 272.08 L1082.46 298.65 L1101.7 317.62 L1136.0699 308.24 L1139.72 294.11 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1601.08 257.8 L1610.75 284.8 L1607.84 291.38 L1569.7 302.94 L1550.95 272.79 L1576.13 252.07 L1601.08 257.8 Z"
      /><path d="M1601.08 257.8 L1610.75 284.8 L1607.84 291.38 L1569.7 302.94 L1550.95 272.79 L1576.13 252.07 L1601.08 257.8 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1142.4 877.99 L1170.33 899.13 L1169.4 917.75 L1133.7 932.8 L1119.51 898.27 L1142.4 877.99 Z"
      /><path d="M1142.4 877.99 L1170.33 899.13 L1169.4 917.75 L1133.7 932.8 L1119.51 898.27 L1142.4 877.99 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M812.13 935.41 L824.35 961.39 L811.46 988.76 L803.52 991.77 L775.3 981.35 L766.93 949.45 L773 939.25 L812.13 935.41 Z"
      /><path d="M812.13 935.41 L824.35 961.39 L811.46 988.76 L803.52 991.77 L775.3 981.35 L766.93 949.45 L773 939.25 L812.13 935.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M681.12 97.42 L689.01 147.67 L674.77 157.64 L638.35 145.03 L642.32 100.73 L681.12 97.42 Z"
      /><path d="M681.12 97.42 L689.01 147.67 L674.77 157.64 L638.35 145.03 L642.32 100.73 L681.12 97.42 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M981.79 972.02 L973.36 970.28 L941.18 993.83 L940.97 996.41 L968.54 1031.25 L982.75 1030.75 L1001.66 1012.65 L981.79 972.02 Z"
      /><path d="M981.79 972.02 L973.36 970.28 L941.18 993.83 L940.97 996.41 L968.54 1031.25 L982.75 1030.75 L1001.66 1012.65 L981.79 972.02 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1741.42 1020.41 L1684.42 1041.64 L1668.58 1021.83 L1677.77 986.89 L1724.85 974.55 L1741.42 1020.41 Z"
      /><path d="M1741.42 1020.41 L1684.42 1041.64 L1668.58 1021.83 L1677.77 986.89 L1724.85 974.55 L1741.42 1020.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M640.93 644.84 L616.99 622.23 L593.45 627.44 L584.23 646.89 L598.66 674.42 L627.19 672.96 L640.93 644.84 Z"
      /><path d="M640.93 644.84 L616.99 622.23 L593.45 627.44 L584.23 646.89 L598.66 674.42 L627.19 672.96 L640.93 644.84 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M363.82 632.41 L340.59 630.61 L325.12 653.07 L347.75 691.29 L377.17 681.08 L384.14 662.38 L363.82 632.41 Z"
      /><path d="M363.82 632.41 L340.59 630.61 L325.12 653.07 L347.75 691.29 L377.17 681.08 L384.14 662.38 L363.82 632.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M950.05 111.25 L930.11 83.67 L905.59 97.05 L907.38 121.6 L937.75 128.48 L950.05 111.25 Z"
      /><path d="M950.05 111.25 L930.11 83.67 L905.59 97.05 L907.38 121.6 L937.75 128.48 L950.05 111.25 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1488.3101 307.47 L1466.98 279.68 L1437.24 283.59 L1432.45 289.08 L1442.35 338.01 L1465.2 341.71 L1488.3101 307.47 Z"
      /><path d="M1488.3101 307.47 L1466.98 279.68 L1437.24 283.59 L1432.45 289.08 L1442.35 338.01 L1465.2 341.71 L1488.3101 307.47 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1221.15 747.73 L1196.42 721.82 L1168.15 731.16 L1162.52 763.16 L1180.92 783.59 L1215.47 776.05 L1221.15 747.73 Z"
      /><path d="M1221.15 747.73 L1196.42 721.82 L1168.15 731.16 L1162.52 763.16 L1180.92 783.59 L1215.47 776.05 L1221.15 747.73 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1600.45 820.23 L1568.92 806.78 L1566 807.77 L1552.8 836.35 L1583.47 868.37 L1601.5 854.96 L1600.45 820.23 Z"
      /><path d="M1600.45 820.23 L1568.92 806.78 L1566 807.77 L1552.8 836.35 L1583.47 868.37 L1601.5 854.96 L1600.45 820.23 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M691.35 928.26 L671.4 904.58 L629.93 919.28 L645.09 952.92 L669.39 959.85 L691.35 928.26 Z"
      /><path d="M691.35 928.26 L671.4 904.58 L629.93 919.28 L645.09 952.92 L669.39 959.85 L691.35 928.26 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M860.07 961.8 L824.35 961.39 L811.46 988.76 L840.3 1008.58 L872.5 990.99 L860.07 961.8 Z"
      /><path d="M860.07 961.8 L824.35 961.39 L811.46 988.76 L840.3 1008.58 L872.5 990.99 L860.07 961.8 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1828.1801 440.17 L1826.74 478.49 L1815.5601 483.61 L1776.02 461.75 L1774.8 446.52 L1810.09 425.14 L1828.1801 440.17 Z"
      /><path d="M1828.1801 440.17 L1826.74 478.49 L1815.5601 483.61 L1776.02 461.75 L1774.8 446.52 L1810.09 425.14 L1828.1801 440.17 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M80.6 363.28 L92.54 374.47 L90.71 414.15 L63.02 421.69 L43.42 401.24 L47.09 371.1 L80.6 363.28 Z"
      /><path d="M80.6 363.28 L92.54 374.47 L90.71 414.15 L63.02 421.69 L43.42 401.24 L47.09 371.1 L80.6 363.28 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1321.41 375.04 L1301.5 413.86 L1301.76 415.95 L1359.45 428.61 L1365.66 422.98 L1368.3 384.07 L1367.0601 382.52 L1321.41 375.04 Z"
      /><path d="M1321.41 375.04 L1301.5 413.86 L1301.76 415.95 L1359.45 428.61 L1365.66 422.98 L1368.3 384.07 L1367.0601 382.52 L1321.41 375.04 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1889.04 306.35 L1878.16 346.08 L1853 350.38 L1844.87 345.48 L1839.52 307.88 L1876.25 296.22 L1889.04 306.35 Z"
      /><path d="M1889.04 306.35 L1878.16 346.08 L1853 350.38 L1844.87 345.48 L1839.52 307.88 L1876.25 296.22 L1889.04 306.35 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M842.95 589.17 L825.12 610.23 L792.98 607.6 L781.64 577.68 L813.79 557.64 L842.95 589.17 Z"
      /><path d="M842.95 589.17 L825.12 610.23 L792.98 607.6 L781.64 577.68 L813.79 557.64 L842.95 589.17 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1578.48 86.3 L1537.76 88.95 L1535.55 122.04 L1572.36 132.14 L1579.45 126.72 L1578.48 86.3 Z"
      /><path d="M1578.48 86.3 L1537.76 88.95 L1535.55 122.04 L1572.36 132.14 L1579.45 126.72 L1578.48 86.3 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M246.97 573.41 L286.91 590.23 L290.51 600.39 L277.53 626.61 L260.22 632.73 L231.39 619.33 L237.33 579.2 L246.97 573.41 Z"
      /><path d="M246.97 573.41 L286.91 590.23 L290.51 600.39 L277.53 626.61 L260.22 632.73 L231.39 619.33 L237.33 579.2 L246.97 573.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M933.02 72.36 L919.69 53.37 L891.85 60.73 L887.69 86.1 L905.59 97.05 L930.11 83.67 L933.02 72.36 Z"
      /><path d="M933.02 72.36 L919.69 53.37 L891.85 60.73 L887.69 86.1 L905.59 97.05 L930.11 83.67 L933.02 72.36 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M70.44 112.18 L76.99 112.21 L100.82 143.49 L98.03 150.45 L63.76 161.34 L58.98 158.75 L55.06 124.7 L70.44 112.18 Z"
      /><path d="M70.44 112.18 L76.99 112.21 L100.82 143.49 L98.03 150.45 L63.76 161.34 L58.98 158.75 L55.06 124.7 L70.44 112.18 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1596.96 677.49 L1577.45 674.82 L1562.88 708.94 L1579.21 727.43 L1601.1801 722.35 L1611.78 695.81 L1596.96 677.49 Z"
      /><path d="M1596.96 677.49 L1577.45 674.82 L1562.88 708.94 L1579.21 727.43 L1601.1801 722.35 L1611.78 695.81 L1596.96 677.49 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M254.08 670.77 L239.36 680.64 L240.68 702.81 L264.03 719.36 L295.2 703.57 L289.8 681.11 L254.08 670.77 Z"
      /><path d="M254.08 670.77 L239.36 680.64 L240.68 702.81 L264.03 719.36 L295.2 703.57 L289.8 681.11 L254.08 670.77 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1236.6801 643.75 L1205.76 641.62 L1185.37 670.21 L1204.77 697.74 L1237.0699 690.06 L1245.66 655.7 L1236.6801 643.75 Z"
      /><path d="M1236.6801 643.75 L1205.76 641.62 L1185.37 670.21 L1204.77 697.74 L1237.0699 690.06 L1245.66 655.7 L1236.6801 643.75 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M527.97 608.02 L540.07 613.4 L549.13 651.42 L540.59 663.3 L523.19 667.27 L495.46 636.55 L502.5 618.66 L527.97 608.02 Z"
      /><path d="M527.97 608.02 L540.07 613.4 L549.13 651.42 L540.59 663.3 L523.19 667.27 L495.46 636.55 L502.5 618.66 L527.97 608.02 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M726.75 198.67 L707.76 211.4 L704.5 242.05 L752.48 261.1 L762.93 247.53 L758.09 212.02 L726.75 198.67 Z"
      /><path d="M726.75 198.67 L707.76 211.4 L704.5 242.05 L752.48 261.1 L762.93 247.53 L758.09 212.02 L726.75 198.67 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M665.55 1028.35 L649.26 1044.41 L654 1080 L690.9 1080 L692.2 1035.17 L665.55 1028.35 Z"
      /><path d="M665.55 1028.35 L649.26 1044.41 L654 1080 L690.9 1080 L692.2 1035.17 L665.55 1028.35 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1014.77 171.79 L985.09 143.44 L959.34 161.09 L962.25 174.19 L990.28 191.51 L1013.26 177.72 L1014.77 171.79 Z"
      /><path d="M1014.77 171.79 L985.09 143.44 L959.34 161.09 L962.25 174.19 L990.28 191.51 L1013.26 177.72 L1014.77 171.79 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1479.9301 255.26 L1448.89 225.56 L1424.98 241.12 L1437.24 283.59 L1466.98 279.68 L1479.9301 255.26 Z"
      /><path d="M1479.9301 255.26 L1448.89 225.56 L1424.98 241.12 L1437.24 283.59 L1466.98 279.68 L1479.9301 255.26 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M278.6 277.5 L251.51 257.39 L231.31 264.78 L234.78 304.04 L262.07 313.98 L278.6 277.5 Z"
      /><path d="M278.6 277.5 L251.51 257.39 L231.31 264.78 L234.78 304.04 L262.07 313.98 L278.6 277.5 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M89.28 763.43 L120.99 777.28 L123.38 815.88 L78.84 831.05 L59.63 808.74 L61.75 776.75 L89.28 763.43 Z"
      /><path d="M89.28 763.43 L120.99 777.28 L123.38 815.88 L78.84 831.05 L59.63 808.74 L61.75 776.75 L89.28 763.43 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M575.69 224.19 L522.29 218.74 L512.13 230.52 L512.95 244.17 L549.14 273.54 L579.02 240.46 L575.69 224.19 Z"
      /><path d="M575.69 224.19 L522.29 218.74 L512.13 230.52 L512.95 244.17 L549.14 273.54 L579.02 240.46 L575.69 224.19 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M289.56 74.7 L309.03 99.61 L305.2 114.94 L275.98 132.95 L252.83 121.47 L248.47 113.3 L253.93 89.53 L289.56 74.7 Z"
      /><path d="M289.56 74.7 L309.03 99.61 L305.2 114.94 L275.98 132.95 L252.83 121.47 L248.47 113.3 L253.93 89.53 L289.56 74.7 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1884.54 576.37 L1920 582.5 L1920 619.5 L1873.03 615.44 L1868.6801 595.2 L1884.54 576.37 Z"
      /><path d="M1884.54 576.37 L1920 582.5 L1920 619.5 L1873.03 615.44 L1868.6801 595.2 L1884.54 576.37 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1442.35 338.01 L1465.2 341.71 L1482.1899 366.03 L1478.49 383.39 L1435.89 408.07 L1416.62 380.45 L1424.74 348.3 L1442.35 338.01 Z"
      /><path d="M1442.35 338.01 L1465.2 341.71 L1482.1899 366.03 L1478.49 383.39 L1435.89 408.07 L1416.62 380.45 L1424.74 348.3 L1442.35 338.01 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1307.52 1023.22 L1333.4 1037.48 L1331.9 1080 L1277.4 1080 L1291.36 1029.33 L1307.52 1023.22 Z"
      /><path d="M1307.52 1023.22 L1333.4 1037.48 L1331.9 1080 L1277.4 1080 L1291.36 1029.33 L1307.52 1023.22 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M216.95 835.55 L213.95 853.95 L183.41 873.91 L147.25 853.53 L144.38 830.79 L178 810.2 L216.95 835.55 Z"
      /><path d="M216.95 835.55 L213.95 853.95 L183.41 873.91 L147.25 853.53 L144.38 830.79 L178 810.2 L216.95 835.55 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1305.42 554.08 L1322.76 566.95 L1325.14 588.32 L1283.09 605.37 L1277.6899 601.94 L1274.72 568.38 L1305.42 554.08 Z"
      /><path d="M1305.42 554.08 L1322.76 566.95 L1325.14 588.32 L1283.09 605.37 L1277.6899 601.94 L1274.72 568.38 L1305.42 554.08 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1387.1 951.67 L1372.8199 987.48 L1420.36 1008.66 L1432.4 994.24 L1430.4399 959.72 L1387.1 951.67 Z"
      /><path d="M1387.1 951.67 L1372.8199 987.48 L1420.36 1008.66 L1432.4 994.24 L1430.4399 959.72 L1387.1 951.67 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1601.11 908.48 L1581.84 873.78 L1548.49 890.21 L1549.3101 924.65 L1576.95 937.25 L1601.11 908.48 Z"
      /><path d="M1601.11 908.48 L1581.84 873.78 L1548.49 890.21 L1549.3101 924.65 L1576.95 937.25 L1601.11 908.48 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M815.8 545.16 L784.17 519.21 L764.23 530.54 L770.77 573.56 L781.64 577.68 L813.79 557.64 L815.8 545.16 Z"
      /><path d="M815.8 545.16 L784.17 519.21 L764.23 530.54 L770.77 573.56 L781.64 577.68 L813.79 557.64 L815.8 545.16 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M240.68 702.81 L264.03 719.36 L262.14 753.6 L255.54 760.6 L209.29 730.02 L240.68 702.81 Z"
      /><path d="M240.68 702.81 L264.03 719.36 L262.14 753.6 L255.54 760.6 L209.29 730.02 L240.68 702.81 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1653 0 L1598 0 L1599.71 40.65 L1640.55 49.3 L1653 0 Z"
      /><path d="M1653 0 L1598 0 L1599.71 40.65 L1640.55 49.3 L1653 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1553.4399 524.47 L1550.25 559.79 L1530.1899 568.93 L1505.87 557.37 L1509.62 522.51 L1544.47 515.82 L1553.4399 524.47 Z"
      /><path d="M1553.4399 524.47 L1550.25 559.79 L1530.1899 568.93 L1505.87 557.37 L1509.62 522.51 L1544.47 515.82 L1553.4399 524.47 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1736.39 621.14 L1747.77 631.46 L1738.15 671.08 L1715.08 669.86 L1700.05 648.99 L1715.5699 622.87 L1736.39 621.14 Z"
      /><path d="M1736.39 621.14 L1747.77 631.46 L1738.15 671.08 L1715.08 669.86 L1700.05 648.99 L1715.5699 622.87 L1736.39 621.14 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M51.3 659.49 L0 659.2 L0 710.2 L43.64 714.75 L51.3 709.24 L51.3 659.49 Z"
      /><path d="M51.3 659.49 L0 659.2 L0 710.2 L43.64 714.75 L51.3 709.24 L51.3 659.49 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M732.37 671.54 L708.41 646.26 L679.28 653.48 L677.35 691.73 L715.15 697.93 L732.37 671.54 Z"
      /><path d="M732.37 671.54 L708.41 646.26 L679.28 653.48 L677.35 691.73 L715.15 697.93 L732.37 671.54 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1419.49 24.85 L1443.75 40.39 L1434.55 71.89 L1395.3 58.58 L1392.8101 48.56 L1419.49 24.85 Z"
      /><path d="M1419.49 24.85 L1443.75 40.39 L1434.55 71.89 L1395.3 58.58 L1392.8101 48.56 L1419.49 24.85 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M91.58 717.52 L51.3 709.24 L43.64 714.75 L42.15 762.81 L61.75 776.75 L89.28 763.43 L91.58 717.52 Z"
      /><path d="M91.58 717.52 L51.3 709.24 L43.64 714.75 L42.15 762.81 L61.75 776.75 L89.28 763.43 L91.58 717.52 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M606.74 852.21 L579.39 862.48 L574.09 878.67 L583.07 897.17 L618.61 902.53 L627.41 869.85 L606.74 852.21 Z"
      /><path d="M606.74 852.21 L579.39 862.48 L574.09 878.67 L583.07 897.17 L618.61 902.53 L627.41 869.85 L606.74 852.21 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1433.5699 482.78 L1438.78 514.74 L1404.45 537.68 L1380.76 501.69 L1386.13 484.95 L1409.78 472.26 L1433.5699 482.78 Z"
      /><path d="M1433.5699 482.78 L1438.78 514.74 L1404.45 537.68 L1380.76 501.69 L1386.13 484.95 L1409.78 472.26 L1433.5699 482.78 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M447.68 310.39 L418.45 287.56 L395.27 299.37 L391.92 313.05 L405.74 337.96 L425.28 339.7 L448.01 312.51 L447.68 310.39 Z"
      /><path d="M447.68 310.39 L418.45 287.56 L395.27 299.37 L391.92 313.05 L405.74 337.96 L425.28 339.7 L448.01 312.51 L447.68 310.39 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M232.91 786.42 L230.73 824.75 L216.95 835.55 L178 810.2 L183.51 774.17 L187.8 771.72 L232.91 786.42 Z"
      /><path d="M232.91 786.42 L230.73 824.75 L216.95 835.55 L178 810.2 L183.51 774.17 L187.8 771.72 L232.91 786.42 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1062.6 0 L1087.9301 40.84 L1119.75 16.6 L1121.2 0 L1062.6 0 Z"
      /><path d="M1062.6 0 L1087.9301 40.84 L1119.75 16.6 L1121.2 0 L1062.6 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M142.69 381.18 L129.93 366.74 L92.54 374.47 L90.71 414.15 L100.48 419.51 L139.94 402.42 L142.69 381.18 Z"
      /><path d="M142.69 381.18 L129.93 366.74 L92.54 374.47 L90.71 414.15 L100.48 419.51 L139.94 402.42 L142.69 381.18 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1323.37 473.87 L1295.8101 428.11 L1275.71 439.44 L1267.51 472.16 L1292.21 490.02 L1323.37 473.87 Z"
      /><path d="M1323.37 473.87 L1295.8101 428.11 L1275.71 439.44 L1267.51 472.16 L1292.21 490.02 L1323.37 473.87 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M870.53 899.39 L863.13 916.03 L820.83 918.6 L810.8 890.77 L828.26 866.42 L845.67 865.35 L870.53 899.39 Z"
      /><path d="M870.53 899.39 L863.13 916.03 L820.83 918.6 L810.8 890.77 L828.26 866.42 L845.67 865.35 L870.53 899.39 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M305.67 336.38 L285.58 371.81 L312.2 390.58 L335.6 377 L335.6 346.82 L305.67 336.38 Z"
      /><path d="M305.67 336.38 L285.58 371.81 L312.2 390.58 L335.6 377 L335.6 346.82 L305.67 336.38 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M446.53 541.53 L438.25 579.34 L450.86 597.03 L477.72 590.95 L491.54 564.82 L486.4 551.71 L446.53 541.53 Z"
      /><path d="M446.53 541.53 L438.25 579.34 L450.86 597.03 L477.72 590.95 L491.54 564.82 L486.4 551.71 L446.53 541.53 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1169.4 917.75 L1187.84 934.68 L1186.78 954.04 L1168.08 968.97 L1141.4399 959.62 L1133.1899 934.15 L1133.7 932.8 L1169.4 917.75 Z"
      /><path d="M1169.4 917.75 L1187.84 934.68 L1186.78 954.04 L1168.08 968.97 L1141.4399 959.62 L1133.1899 934.15 L1133.7 932.8 L1169.4 917.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M726.71 813.38 L754.18 816.75 L768.11 851.21 L766.24 855.73 L714.68 866.34 L713.54 865.6 L708.1 839.98 L726.71 813.38 Z"
      /><path d="M726.71 813.38 L754.18 816.75 L768.11 851.21 L766.24 855.73 L714.68 866.34 L713.54 865.6 L708.1 839.98 L726.71 813.38 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M115.71 1030.67 L92.85 991.55 L61.1 992.87 L50.77 1012.27 L57.47 1043.63 L57.54 1043.71 L113.78 1034.2 L115.71 1030.67 Z"
      /><path d="M115.71 1030.67 L92.85 991.55 L61.1 992.87 L50.77 1012.27 L57.47 1043.63 L57.54 1043.71 L113.78 1034.2 L115.71 1030.67 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1267.51 472.16 L1292.21 490.02 L1289.8199 515.82 L1263.67 525.19 L1242.08 509.3 L1245.58 480.74 L1267.51 472.16 Z"
      /><path d="M1267.51 472.16 L1292.21 490.02 L1289.8199 515.82 L1263.67 525.19 L1242.08 509.3 L1245.58 480.74 L1267.51 472.16 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1222.4399 364.42 L1246.5601 381.9 L1232.65 422.34 L1224.53 427.21 L1195.22 418.54 L1182.08 386.85 L1187.45 375.94 L1222.4399 364.42 Z"
      /><path d="M1222.4399 364.42 L1246.5601 381.9 L1232.65 422.34 L1224.53 427.21 L1195.22 418.54 L1182.08 386.85 L1187.45 375.94 L1222.4399 364.42 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M718.37 614.82 L692.88 597.46 L669.86 606.61 L661.97 640.38 L679.28 653.48 L708.41 646.26 L718.37 614.82 Z"
      /><path d="M718.37 614.82 L692.88 597.46 L669.86 606.61 L661.97 640.38 L679.28 653.48 L708.41 646.26 L718.37 614.82 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1221.03 181.57 L1205.48 143.66 L1177.91 146.08 L1167.9 164.4 L1183.08 194.23 L1216.65 188.6 L1221.03 181.57 Z"
      /><path d="M1221.03 181.57 L1205.48 143.66 L1177.91 146.08 L1167.9 164.4 L1183.08 194.23 L1216.65 188.6 L1221.03 181.57 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M110.36 177.97 L130.63 181.81 L139 210.26 L109.45 229.29 L92.46 196.84 L110.36 177.97 Z"
      /><path d="M110.36 177.97 L130.63 181.81 L139 210.26 L109.45 229.29 L92.46 196.84 L110.36 177.97 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M385.1 362.8 L385.14 368.51 L360.13 389.86 L335.6 377 L335.6 346.82 L351.99 336.07 L385.1 362.8 Z"
      /><path d="M385.1 362.8 L385.14 368.51 L360.13 389.86 L335.6 377 L335.6 346.82 L351.99 336.07 L385.1 362.8 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M470.92 712.95 L494.57 738.83 L492.8 754.37 L455.54 767.65 L439.41 752.39 L446.42 718.75 L470.92 712.95 Z"
      /><path d="M470.92 712.95 L494.57 738.83 L492.8 754.37 L455.54 767.65 L439.41 752.39 L446.42 718.75 L470.92 712.95 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M770.77 573.56 L746.56 582.18 L735.31 609.58 L766.62 634.9 L775.54 633.3 L792.98 607.6 L781.64 577.68 L770.77 573.56 Z"
      /><path d="M770.77 573.56 L746.56 582.18 L735.31 609.58 L766.62 634.9 L775.54 633.3 L792.98 607.6 L781.64 577.68 L770.77 573.56 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1445.65 737.03 L1433.46 760.75 L1413.1801 760.19 L1396.21 737.57 L1408.5601 710.98 L1428.8 708.05 L1445.65 737.03 Z"
      /><path d="M1445.65 737.03 L1433.46 760.75 L1413.1801 760.19 L1396.21 737.57 L1408.5601 710.98 L1428.8 708.05 L1445.65 737.03 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1183.55 849 L1143.17 861.32 L1142.4 877.99 L1170.33 899.13 L1196.05 880.8 L1183.55 849 Z"
      /><path d="M1183.55 849 L1143.17 861.32 L1142.4 877.99 L1170.33 899.13 L1196.05 880.8 L1183.55 849 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1182.08 386.85 L1195.22 418.54 L1166.01 446.57 L1136.02 424.95 L1145 393.03 L1182.08 386.85 Z"
      /><path d="M1182.08 386.85 L1195.22 418.54 L1166.01 446.57 L1136.02 424.95 L1145 393.03 L1182.08 386.85 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M362.87 413.88 L378.52 423 L383.32 456.18 L370.85 468.92 L335.35 463.79 L335.43 429.57 L362.87 413.88 Z"
      /><path d="M362.87 413.88 L378.52 423 L383.32 456.18 L370.85 468.92 L335.35 463.79 L335.43 429.57 L362.87 413.88 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M301.79 990.77 L338.31 1008.3 L339.26 1030.47 L319.62 1049.8199 L282.63 1030.8199 L281.63 1007.9 L301.79 990.77 Z"
      /><path d="M301.79 990.77 L338.31 1008.3 L339.26 1030.47 L319.62 1049.8199 L282.63 1030.8199 L281.63 1007.9 L301.79 990.77 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M149.63 603.43 L124.92 627.38 L103.2 624.55 L86.79 590.7 L95.5 576.8 L135.95 570.82 L149.63 603.43 Z"
      /><path d="M149.63 603.43 L124.92 627.38 L103.2 624.55 L86.79 590.7 L95.5 576.8 L135.95 570.82 L149.63 603.43 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M858.21 485.7 L835.42 501.16 L836.94 529.63 L869.15 542.3 L887.61 501.45 L858.21 485.7 Z"
      /><path d="M858.21 485.7 L835.42 501.16 L836.94 529.63 L869.15 542.3 L887.61 501.45 L858.21 485.7 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M393.92 579.01 L438.25 579.34 L450.86 597.03 L444.97 614.6 L419.65 627.06 L389.85 604.2 L388.46 584.77 L393.92 579.01 Z"
      /><path d="M393.92 579.01 L438.25 579.34 L450.86 597.03 L444.97 614.6 L419.65 627.06 L389.85 604.2 L388.46 584.77 L393.92 579.01 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M523.98 572.82 L491.54 564.82 L477.72 590.95 L502.5 618.66 L527.97 608.02 L523.98 572.82 Z"
      /><path d="M523.98 572.82 L491.54 564.82 L477.72 590.95 L502.5 618.66 L527.97 608.02 L523.98 572.82 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M613.74 1037.5699 L649.26 1044.41 L654 1080 L606.3 1080 L613.74 1037.5699 Z"
      /><path d="M613.74 1037.5699 L649.26 1044.41 L654 1080 L606.3 1080 L613.74 1037.5699 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M996.81 691 L1047.13 701.58 L1049.04 704.4 L1046.26 723.17 L1014.68 747.47 L999 744.52 L988.16 727.94 L996.81 691 Z"
      /><path d="M996.81 691 L1047.13 701.58 L1049.04 704.4 L1046.26 723.17 L1014.68 747.47 L999 744.52 L988.16 727.94 L996.81 691 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M526.15 301.36 L504.94 301.01 L487.96 332.19 L520.45 351.88 L543.75 336.54 L526.15 301.36 Z"
      /><path d="M526.15 301.36 L504.94 301.01 L487.96 332.19 L520.45 351.88 L543.75 336.54 L526.15 301.36 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M342.87 298.13 L326.64 291.37 L317.91 294.11 L301.57 327.21 L305.67 336.38 L335.6 346.82 L351.99 336.07 L355.09 325.55 L342.87 298.13 Z"
      /><path d="M342.87 298.13 L326.64 291.37 L317.91 294.11 L301.57 327.21 L305.67 336.38 L335.6 346.82 L351.99 336.07 L355.09 325.55 L342.87 298.13 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1725.12 219.18 L1742.04 222.3 L1755.76 250.33 L1736.47 270.39 L1705.99 265.71 L1697.9 243.59 L1725.12 219.18 Z"
      /><path d="M1725.12 219.18 L1742.04 222.3 L1755.76 250.33 L1736.47 270.39 L1705.99 265.71 L1697.9 243.59 L1725.12 219.18 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M377.17 681.08 L401.54 708.16 L390.45 735.12 L359.56 738.1 L342.34 701.86 L347.75 691.29 L377.17 681.08 Z"
      /><path d="M377.17 681.08 L401.54 708.16 L390.45 735.12 L359.56 738.1 L342.34 701.86 L347.75 691.29 L377.17 681.08 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1616.85 443.42 L1580.14 432.67 L1573.34 437.05 L1565.23 469.67 L1598.05 491.93 L1623.87 482.73 L1624.72 481.14 L1616.85 443.42 Z"
      /><path d="M1616.85 443.42 L1580.14 432.67 L1573.34 437.05 L1565.23 469.67 L1598.05 491.93 L1623.87 482.73 L1624.72 481.14 L1616.85 443.42 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M766.62 634.9 L735.31 609.58 L718.37 614.82 L708.41 646.26 L732.37 671.54 L745.96 669.76 L766.62 634.9 Z"
      /><path d="M766.62 634.9 L735.31 609.58 L718.37 614.82 L708.41 646.26 L732.37 671.54 L745.96 669.76 L766.62 634.9 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M826.61 806.98 L850.42 810.78 L864.87 842.26 L845.67 865.35 L828.26 866.42 L807.25 836.89 L812.16 818.03 L826.61 806.98 Z"
      /><path d="M826.61 806.98 L850.42 810.78 L864.87 842.26 L845.67 865.35 L828.26 866.42 L807.25 836.89 L812.16 818.03 L826.61 806.98 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1062.6 0 L1054.4 0 L1035.88 37.08 L1040.23 50.28 L1063.12 62.24 L1086.89 48.06 L1087.9301 40.84 L1062.6 0 Z"
      /><path d="M1062.6 0 L1054.4 0 L1035.88 37.08 L1040.23 50.28 L1063.12 62.24 L1086.89 48.06 L1087.9301 40.84 L1062.6 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1529.3199 80.05 L1495.9399 87.72 L1488.72 115.82 L1492.3101 121.4 L1524.22 131.58 L1535.55 122.04 L1537.76 88.95 L1529.3199 80.05 Z"
      /><path d="M1529.3199 80.05 L1495.9399 87.72 L1488.72 115.82 L1492.3101 121.4 L1524.22 131.58 L1535.55 122.04 L1537.76 88.95 L1529.3199 80.05 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1122.88 147.29 L1137.1801 168.66 L1127.17 196.34 L1117.75 201.94 L1080.6801 173.93 L1092.24 149.06 L1122.88 147.29 Z"
      /><path d="M1122.88 147.29 L1137.1801 168.66 L1127.17 196.34 L1117.75 201.94 L1080.6801 173.93 L1092.24 149.06 L1122.88 147.29 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1741.42 1020.41 L1750.85 1025.92 L1753.5 1080 L1684.1 1080 L1684.42 1041.64 L1741.42 1020.41 Z"
      /><path d="M1741.42 1020.41 L1750.85 1025.92 L1753.5 1080 L1684.1 1080 L1684.42 1041.64 L1741.42 1020.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M217.6 490.94 L227.9 518.33 L191.45 545.43 L164.76 495.83 L165.34 493.73 L173.17 487.85 L217.6 490.94 Z"
      /><path d="M217.6 490.94 L227.9 518.33 L191.45 545.43 L164.76 495.83 L165.34 493.73 L173.17 487.85 L217.6 490.94 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M549.36 553.89 L546.29 553.73 L523.98 572.82 L527.97 608.02 L540.07 613.4 L571.96 599.49 L575.72 585.44 L549.36 553.89 Z"
      /><path d="M549.36 553.89 L546.29 553.73 L523.98 572.82 L527.97 608.02 L540.07 613.4 L571.96 599.49 L575.72 585.44 L549.36 553.89 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 242.1 L1920 178 L1883.54 184.29 L1871.84 207.17 L1920 242.1 Z"
      /><path d="M1920 242.1 L1920 178 L1883.54 184.29 L1871.84 207.17 L1920 242.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1478.36 159.64 L1454.28 158.16 L1438.21 188.04 L1453.1801 209.61 L1481.5 201.87 L1492.88 174.36 L1478.36 159.64 Z"
      /><path d="M1478.36 159.64 L1454.28 158.16 L1438.21 188.04 L1453.1801 209.61 L1481.5 201.87 L1492.88 174.36 L1478.36 159.64 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M470.77 646.38 L463.86 663.1 L434.33 670.95 L414.83 652.42 L419.65 627.06 L444.97 614.6 L470.77 646.38 Z"
      /><path d="M470.77 646.38 L463.86 663.1 L434.33 670.95 L414.83 652.42 L419.65 627.06 L444.97 614.6 L470.77 646.38 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M477.72 590.95 L450.86 597.03 L444.97 614.6 L470.77 646.38 L495.46 636.55 L502.5 618.66 L477.72 590.95 Z"
      /><path d="M477.72 590.95 L450.86 597.03 L444.97 614.6 L470.77 646.38 L495.46 636.55 L502.5 618.66 L477.72 590.95 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M891.65 146.96 L916.46 167.32 L913.66 187.04 L887.48 198.28 L875.55 191.79 L869.9 161.34 L891.65 146.96 Z"
      /><path d="M891.65 146.96 L916.46 167.32 L913.66 187.04 L887.48 198.28 L875.55 191.79 L869.9 161.34 L891.65 146.96 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1166.01 446.57 L1168.1899 467.78 L1149.99 483.05 L1117 478.95 L1103.6899 456.55 L1111.52 433.34 L1136.02 424.95 L1166.01 446.57 Z"
      /><path d="M1166.01 446.57 L1168.1899 467.78 L1149.99 483.05 L1117 478.95 L1103.6899 456.55 L1111.52 433.34 L1136.02 424.95 L1166.01 446.57 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1792.24 976.03 L1775.95 952.44 L1725.75 972.5 L1724.85 974.55 L1741.42 1020.41 L1750.85 1025.92 L1776.91 1017.54 L1792.24 976.03 Z"
      /><path d="M1792.24 976.03 L1775.95 952.44 L1725.75 972.5 L1724.85 974.55 L1741.42 1020.41 L1750.85 1025.92 L1776.91 1017.54 L1792.24 976.03 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M468.84 449.46 L453.87 424.48 L427.16 428.26 L415.99 459.54 L426.41 474.82 L448.8 475.17 L468.84 449.46 Z"
      /><path d="M468.84 449.46 L453.87 424.48 L427.16 428.26 L415.99 459.54 L426.41 474.82 L448.8 475.17 L468.84 449.46 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M367.78 832.42 L354.92 810.43 L323.56 814.24 L314.76 849.93 L337.43 869.88 L345.55 869.3 L367.78 832.42 Z"
      /><path d="M367.78 832.42 L354.92 810.43 L323.56 814.24 L314.76 849.93 L337.43 869.88 L345.55 869.3 L367.78 832.42 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M714.68 866.34 L728.43 904.21 L710.43 928.48 L691.35 928.26 L671.4 904.58 L674.67 881.7 L713.54 865.6 L714.68 866.34 Z"
      /><path d="M714.68 866.34 L728.43 904.21 L710.43 928.48 L691.35 928.26 L671.4 904.58 L674.67 881.7 L713.54 865.6 L714.68 866.34 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1530.1899 568.93 L1505.87 557.37 L1492.04 564.03 L1488.24 611.46 L1488.85 612.37 L1495.33 614.46 L1529.54 602.54 L1530.1899 568.93 Z"
      /><path d="M1530.1899 568.93 L1505.87 557.37 L1492.04 564.03 L1488.24 611.46 L1488.85 612.37 L1495.33 614.46 L1529.54 602.54 L1530.1899 568.93 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1072.5601 985.78 L1042.24 976.05 L1020.45 1013.34 L1036.8101 1031.1899 L1057.84 1032.58 L1076.9301 1005.25 L1072.5601 985.78 Z"
      /><path d="M1072.5601 985.78 L1042.24 976.05 L1020.45 1013.34 L1036.8101 1031.1899 L1057.84 1032.58 L1076.9301 1005.25 L1072.5601 985.78 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1121.2 0 L1165.6 0 L1167.66 33.83 L1142.02 45.85 L1119.75 16.6 L1121.2 0 Z"
      /><path d="M1121.2 0 L1165.6 0 L1167.66 33.83 L1142.02 45.85 L1119.75 16.6 L1121.2 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1338.7 0 L1375.6 0 L1377.05 37.54 L1341.35 47.64 L1334.9301 39.94 L1338.7 0 Z"
      /><path d="M1338.7 0 L1375.6 0 L1377.05 37.54 L1341.35 47.64 L1334.9301 39.94 L1338.7 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1336.8101 668.87 L1337.3101 669.32 L1344.97 703.61 L1311.9 720.43 L1287.9301 700.2 L1293.39 675.43 L1336.8101 668.87 Z"
      /><path d="M1336.8101 668.87 L1337.3101 669.32 L1344.97 703.61 L1311.9 720.43 L1287.9301 700.2 L1293.39 675.43 L1336.8101 668.87 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M671.18 799.59 L640.56 769.98 L617.67 783.67 L616.16 816.42 L660.31 827.04 L666.53 822.38 L671.18 799.59 Z"
      /><path d="M671.18 799.59 L640.56 769.98 L617.67 783.67 L616.16 816.42 L660.31 827.04 L666.53 822.38 L671.18 799.59 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M887.69 86.1 L867.87 93.68 L861.92 111.23 L893.5 134.16 L907.38 121.6 L905.59 97.05 L887.69 86.1 Z"
      /><path d="M887.69 86.1 L867.87 93.68 L861.92 111.23 L893.5 134.16 L907.38 121.6 L905.59 97.05 L887.69 86.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1488.4 763.71 L1502.21 798.77 L1471.88 812.56 L1447.8 788.39 L1448.1899 780.85 L1488.4 763.71 Z"
      /><path d="M1488.4 763.71 L1502.21 798.77 L1471.88 812.56 L1447.8 788.39 L1448.1899 780.85 L1488.4 763.71 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M872.35 939.1 L863.13 916.03 L820.83 918.6 L812.13 935.41 L824.35 961.39 L860.07 961.8 L872.35 939.1 Z"
      /><path d="M872.35 939.1 L863.13 916.03 L820.83 918.6 L812.13 935.41 L824.35 961.39 L860.07 961.8 L872.35 939.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1730.49 49.14 L1746.4 89.11 L1740.98 103.56 L1739.89 104.52 L1691.84 92.85 L1684.61 63.43 L1695.16 51.68 L1730.49 49.14 Z"
      /><path d="M1730.49 49.14 L1746.4 89.11 L1740.98 103.56 L1739.89 104.52 L1691.84 92.85 L1684.61 63.43 L1695.16 51.68 L1730.49 49.14 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1537.74 219.4 L1531 214.44 L1502.23 223.75 L1492.97 250.46 L1528.02 271.86 L1535.54 269.29 L1537.74 219.4 Z"
      /><path d="M1537.74 219.4 L1531 214.44 L1502.23 223.75 L1492.97 250.46 L1528.02 271.86 L1535.54 269.29 L1537.74 219.4 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1211.52 21.38 L1180.3199 40.3 L1188.74 62.03 L1234.0601 58.59 L1235.37 55.6 L1211.52 21.38 Z"
      /><path d="M1211.52 21.38 L1180.3199 40.3 L1188.74 62.03 L1234.0601 58.59 L1235.37 55.6 L1211.52 21.38 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M311.67 414.39 L335.43 429.57 L335.35 463.79 L328.89 469.16 L282.39 453.74 L282.77 431.58 L311.67 414.39 Z"
      /><path d="M311.67 414.39 L335.43 429.57 L335.35 463.79 L328.89 469.16 L282.39 453.74 L282.77 431.58 L311.67 414.39 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M33.96 120.8 L13.63 138.41 L37.2 164.54 L58.98 158.75 L55.06 124.7 L33.96 120.8 Z"
      /><path d="M33.96 120.8 L13.63 138.41 L37.2 164.54 L58.98 158.75 L55.06 124.7 L33.96 120.8 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M648.81 42.16 L642.61 46.45 L634.78 93.96 L642.32 100.73 L681.12 97.42 L683.79 94.77 L681.36 52.39 L648.81 42.16 Z"
      /><path d="M648.81 42.16 L642.61 46.45 L634.78 93.96 L642.32 100.73 L681.12 97.42 L683.79 94.77 L681.36 52.39 L648.81 42.16 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1646.73 59.3 L1684.61 63.43 L1691.84 92.85 L1672.52 121.11 L1631.48 99.71 L1630.3101 95.66 L1646.73 59.3 Z"
      /><path d="M1646.73 59.3 L1684.61 63.43 L1691.84 92.85 L1672.52 121.11 L1631.48 99.71 L1630.3101 95.66 L1646.73 59.3 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M820.74 773.07 L785.78 764.01 L772.3 775.8 L772.5 795.16 L812.16 818.03 L826.61 806.98 L820.74 773.07 Z"
      /><path d="M820.74 773.07 L785.78 764.01 L772.3 775.8 L772.5 795.16 L812.16 818.03 L826.61 806.98 L820.74 773.07 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1391.61 858.61 L1383.88 882.02 L1351.87 893.48 L1324.15 871.89 L1331.6 849.42 L1361.03 836.66 L1391.61 858.61 Z"
      /><path d="M1391.61 858.61 L1383.88 882.02 L1351.87 893.48 L1324.15 871.89 L1331.6 849.42 L1361.03 836.66 L1391.61 858.61 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1570.73 751.87 L1584.99 770.94 L1568.92 806.78 L1566 807.77 L1535.9301 789.34 L1538.6899 757.67 L1570.73 751.87 Z"
      /><path d="M1570.73 751.87 L1584.99 770.94 L1568.92 806.78 L1566 807.77 L1535.9301 789.34 L1538.6899 757.67 L1570.73 751.87 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M38.53 333.85 L35.38 359.87 L0 363.9 L0 315.1 L16.16 314.53 L38.53 333.85 Z"
      /><path d="M38.53 333.85 L35.38 359.87 L0 363.9 L0 315.1 L16.16 314.53 L38.53 333.85 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1510.1 802.19 L1502.21 798.77 L1471.88 812.56 L1466.95 836.74 L1485.6801 850.72 L1517.55 836.36 L1510.1 802.19 Z"
      /><path d="M1510.1 802.19 L1502.21 798.77 L1471.88 812.56 L1466.95 836.74 L1485.6801 850.72 L1517.55 836.36 L1510.1 802.19 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1478.49 383.39 L1511.87 423.4 L1464.64 445.41 L1435.39 412.23 L1435.89 408.07 L1478.49 383.39 Z"
      /><path d="M1478.49 383.39 L1511.87 423.4 L1464.64 445.41 L1435.39 412.23 L1435.89 408.07 L1478.49 383.39 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M425.63 928.74 L453.37 930.28 L469.39 952.48 L469.09 955.65 L432.78 984.26 L421.14 981.81 L409.87 960.75 L425.63 928.74 Z"
      /><path d="M425.63 928.74 L453.37 930.28 L469.39 952.48 L469.09 955.65 L432.78 984.26 L421.14 981.81 L409.87 960.75 L425.63 928.74 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1612.27 1003.45 L1557.6 1005.65 L1552.96 1018.15 L1597.6 1080 L1601.6 1080 L1625.95 1023.34 L1612.27 1003.45 Z"
      /><path d="M1612.27 1003.45 L1557.6 1005.65 L1552.96 1018.15 L1597.6 1080 L1601.6 1080 L1625.95 1023.34 L1612.27 1003.45 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M733.4 55.09 L721.06 94.31 L683.79 94.77 L681.36 52.39 L698.26 41.61 L733.4 55.09 Z"
      /><path d="M733.4 55.09 L721.06 94.31 L683.79 94.77 L681.36 52.39 L698.26 41.61 L733.4 55.09 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M996.81 691 L988.16 727.94 L944.27 727.43 L937.27 703.97 L949.66 684.81 L991.48 681.3 L996.81 691 Z"
      /><path d="M996.81 691 L988.16 727.94 L944.27 727.43 L937.27 703.97 L949.66 684.81 L991.48 681.3 L996.81 691 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1107.9301 734.61 L1105.23 743.89 L1074 756.27 L1046.26 723.17 L1049.04 704.4 L1090.24 701.39 L1107.9301 734.61 Z"
      /><path d="M1107.9301 734.61 L1105.23 743.89 L1074 756.27 L1046.26 723.17 L1049.04 704.4 L1090.24 701.39 L1107.9301 734.61 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M936.75 217.86 L951.94 254.88 L941.73 271.16 L904.99 256.18 L901.21 238.61 L936.75 217.86 Z"
      /><path d="M936.75 217.86 L951.94 254.88 L941.73 271.16 L904.99 256.18 L901.21 238.61 L936.75 217.86 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1491.51 980.97 L1472.98 951.28 L1435.6899 954.1 L1430.4399 959.72 L1432.4 994.24 L1482.92 999.72 L1491.51 980.97 Z"
      /><path d="M1491.51 980.97 L1472.98 951.28 L1435.6899 954.1 L1430.4399 959.72 L1432.4 994.24 L1482.92 999.72 L1491.51 980.97 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M691.35 928.26 L710.43 928.48 L727.4 954.25 L717.95 983.19 L708.99 987.94 L676.72 978.29 L669.39 959.85 L691.35 928.26 Z"
      /><path d="M691.35 928.26 L710.43 928.48 L727.4 954.25 L717.95 983.19 L708.99 987.94 L676.72 978.29 L669.39 959.85 L691.35 928.26 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M335.66 150.99 L372.08 175.33 L371.14 197.3 L356.34 208.67 L332.76 206.54 L316.01 187.35 L317.62 169.04 L334.9 151.1 L335.66 150.99 Z"
      /><path d="M335.66 150.99 L372.08 175.33 L371.14 197.3 L356.34 208.67 L332.76 206.54 L316.01 187.35 L317.62 169.04 L334.9 151.1 L335.66 150.99 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M40.69 205.45 L25.48 227.98 L0 229.4 L0 186.2 L26.16 184.86 L40.69 205.45 Z"
      /><path d="M40.69 205.45 L25.48 227.98 L0 229.4 L0 186.2 L26.16 184.86 L40.69 205.45 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M589.47 105.36 L554.16 93.59 L534.98 104.74 L533.77 128.71 L564.85 154.91 L589.86 140.28 L589.47 105.36 Z"
      /><path d="M589.47 105.36 L554.16 93.59 L534.98 104.74 L533.77 128.71 L564.85 154.91 L589.86 140.28 L589.47 105.36 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M812.34 1044.52 L793.69 1031.5 L772.72 1036.89 L769.3 1080 L810.6 1080 L812.34 1044.52 Z"
      /><path d="M812.34 1044.52 L793.69 1031.5 L772.72 1036.89 L769.3 1080 L810.6 1080 L812.34 1044.52 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1669.97 735.46 L1650.48 725.5 L1624.79 742.97 L1623.71 761.78 L1664.47 776.24 L1676 762.72 L1669.97 735.46 Z"
      /><path d="M1669.97 735.46 L1650.48 725.5 L1624.79 742.97 L1623.71 761.78 L1664.47 776.24 L1676 762.72 L1669.97 735.46 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M610.85 821.19 L564.3 812.76 L560.34 838.95 L579.39 862.48 L606.74 852.21 L610.85 821.19 Z"
      /><path d="M610.85 821.19 L564.3 812.76 L560.34 838.95 L579.39 862.48 L606.74 852.21 L610.85 821.19 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 698.2 L1920 652.9 L1872.83 657.57 L1867.6 670.91 L1884.73 700.3 L1920 698.2 Z"
      /><path d="M1920 698.2 L1920 652.9 L1872.83 657.57 L1867.6 670.91 L1884.73 700.3 L1920 698.2 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1321.9 218.59 L1299.6 236.39 L1297.21 266.75 L1300.01 269.75 L1350.8 270.86 L1353.52 268.67 L1345.09 222.99 L1321.9 218.59 Z"
      /><path d="M1321.9 218.59 L1299.6 236.39 L1297.21 266.75 L1300.01 269.75 L1350.8 270.86 L1353.52 268.67 L1345.09 222.99 L1321.9 218.59 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1275.71 439.44 L1232.65 422.34 L1224.53 427.21 L1222.38 464.89 L1245.58 480.74 L1267.51 472.16 L1275.71 439.44 Z"
      /><path d="M1275.71 439.44 L1232.65 422.34 L1224.53 427.21 L1222.38 464.89 L1245.58 480.74 L1267.51 472.16 L1275.71 439.44 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M575.53 370.92 L601.49 390.81 L603.61 419.04 L571.04 434.9 L553.34 428.25 L549.6 393.46 L575.53 370.92 Z"
      /><path d="M575.53 370.92 L601.49 390.81 L603.61 419.04 L571.04 434.9 L553.34 428.25 L549.6 393.46 L575.53 370.92 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1201.15 519.65 L1172.95 535.64 L1173.71 558.86 L1213.5 583.27 L1217.8199 582.09 L1229.52 563.84 L1213.3199 523.34 L1201.15 519.65 Z"
      /><path d="M1201.15 519.65 L1172.95 535.64 L1173.71 558.86 L1213.5 583.27 L1217.8199 582.09 L1229.52 563.84 L1213.3199 523.34 L1201.15 519.65 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M372.15 919.63 L370.22 918.07 L330.59 926.39 L326.25 951.16 L359.87 974.15 L379.2 954.88 L372.15 919.63 Z"
      /><path d="M372.15 919.63 L370.22 918.07 L330.59 926.39 L326.25 951.16 L359.87 974.15 L379.2 954.88 L372.15 919.63 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1706.4301 541.91 L1678.39 536.82 L1660.86 568.85 L1662.66 573.54 L1694.01 590.7 L1712.83 573.46 L1706.4301 541.91 Z"
      /><path d="M1706.4301 541.91 L1678.39 536.82 L1660.86 568.85 L1662.66 573.54 L1694.01 590.7 L1712.83 573.46 L1706.4301 541.91 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1898.47 362.06 L1878.16 346.08 L1853 350.38 L1853 391.78 L1869.71 405.13 L1874.17 403.56 L1898.47 362.06 Z"
      /><path d="M1898.47 362.06 L1878.16 346.08 L1853 350.38 L1853 391.78 L1869.71 405.13 L1874.17 403.56 L1898.47 362.06 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M811.74 455.03 L786.23 442.63 L765.86 451.7 L759.85 474.33 L789.56 498.82 L808.72 488.38 L811.74 455.03 Z"
      /><path d="M811.74 455.03 L786.23 442.63 L765.86 451.7 L759.85 474.33 L789.56 498.82 L808.72 488.38 L811.74 455.03 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M74.19 876.57 L81 881.65 L85.83 935.56 L51.16 949.59 L29.07 914.03 L74.19 876.57 Z"
      /><path d="M74.19 876.57 L81 881.65 L85.83 935.56 L51.16 949.59 L29.07 914.03 L74.19 876.57 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M832.42 199.33 L808.04 212.43 L805.24 244.96 L813.29 253.07 L848.78 250.57 L854.45 240.71 L845.03 205.61 L832.42 199.33 Z"
      /><path d="M832.42 199.33 L808.04 212.43 L805.24 244.96 L813.29 253.07 L848.78 250.57 L854.45 240.71 L845.03 205.61 L832.42 199.33 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M550.9 0 L505.4 0 L504.72 43.19 L513.88 50.08 L548.83 44.72 L550.9 0 Z"
      /><path d="M550.9 0 L505.4 0 L504.72 43.19 L513.88 50.08 L548.83 44.72 L550.9 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1438.21 188.04 L1412.03 185.89 L1393.8199 217.74 L1403.2 235.67 L1424.98 241.12 L1448.89 225.56 L1453.1801 209.61 L1438.21 188.04 Z"
      /><path d="M1438.21 188.04 L1412.03 185.89 L1393.8199 217.74 L1403.2 235.67 L1424.98 241.12 L1448.89 225.56 L1453.1801 209.61 L1438.21 188.04 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1352.8101 547.97 L1369.59 557.15 L1370.8101 585.77 L1336.17 598.08 L1325.14 588.32 L1322.76 566.95 L1352.8101 547.97 Z"
      /><path d="M1352.8101 547.97 L1369.59 557.15 L1370.8101 585.77 L1336.17 598.08 L1325.14 588.32 L1322.76 566.95 L1352.8101 547.97 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M275.64 869.04 L242.61 882.45 L237.46 906.55 L270.79 931.66 L297.27 905.55 L275.64 869.04 Z"
      /><path d="M275.64 869.04 L242.61 882.45 L237.46 906.55 L270.79 931.66 L297.27 905.55 L275.64 869.04 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M25.48 227.98 L0 229.4 L0 267.8 L30.71 271.2 L44.7 253.81 L25.48 227.98 Z"
      /><path d="M25.48 227.98 L0 229.4 L0 267.8 L30.71 271.2 L44.7 253.81 L25.48 227.98 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M939.74 209.75 L913.66 187.04 L887.48 198.28 L891.19 231.55 L901.21 238.61 L936.75 217.86 L939.74 209.75 Z"
      /><path d="M939.74 209.75 L913.66 187.04 L887.48 198.28 L891.19 231.55 L901.21 238.61 L936.75 217.86 L939.74 209.75 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M533.77 128.71 L564.85 154.91 L561.03 171.49 L523.42 187.06 L499.24 166.04 L499.05 151.69 L533.77 128.71 Z"
      /><path d="M533.77 128.71 L564.85 154.91 L561.03 171.49 L523.42 187.06 L499.24 166.04 L499.05 151.69 L533.77 128.71 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1044.47 128.92 L1081.42 130.1 L1092.24 149.06 L1080.6801 173.93 L1070.17 178.46 L1035.97 154.78 L1038 136.43 L1044.47 128.92 Z"
      /><path d="M1044.47 128.92 L1081.42 130.1 L1092.24 149.06 L1080.6801 173.93 L1070.17 178.46 L1035.97 154.78 L1038 136.43 L1044.47 128.92 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M171.68 131.44 L196.81 135.13 L207.23 156.78 L178.73 181.27 L151.11 162.7 L150.72 153.18 L171.68 131.44 Z"
      /><path d="M171.68 131.44 L196.81 135.13 L207.23 156.78 L178.73 181.27 L151.11 162.7 L150.72 153.18 L171.68 131.44 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M878.6 993.78 L872.5 990.99 L840.3 1008.58 L839.72 1034.54 L854.99 1045.95 L875.24 1040.15 L887.54 1012.41 L878.6 993.78 Z"
      /><path d="M878.6 993.78 L872.5 990.99 L840.3 1008.58 L839.72 1034.54 L854.99 1045.95 L875.24 1040.15 L887.54 1012.41 L878.6 993.78 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M302.66 545.21 L255.42 535.85 L246.97 573.41 L286.91 590.23 L306.5 552.95 L302.66 545.21 Z"
      /><path d="M302.66 545.21 L255.42 535.85 L246.97 573.41 L286.91 590.23 L306.5 552.95 L302.66 545.21 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M548.83 44.72 L513.88 50.08 L511.79 90.52 L534.98 104.74 L554.16 93.59 L558.26 52.58 L548.83 44.72 Z"
      /><path d="M548.83 44.72 L513.88 50.08 L511.79 90.52 L534.98 104.74 L554.16 93.59 L558.26 52.58 L548.83 44.72 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M265.5 187.6 L288.99 201.16 L288.56 228.92 L259.4 235.26 L245.91 214.63 L265.5 187.6 Z"
      /><path d="M265.5 187.6 L288.99 201.16 L288.56 228.92 L259.4 235.26 L245.91 214.63 L265.5 187.6 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M529.74 907.42 L512.72 915.98 L509.13 932.56 L527.88 959.67 L551.47 959.1 L568.86 936.52 L566.49 927.27 L529.74 907.42 Z"
      /><path d="M529.74 907.42 L512.72 915.98 L509.13 932.56 L527.88 959.67 L551.47 959.1 L568.86 936.52 L566.49 927.27 L529.74 907.42 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M144.38 830.79 L147.25 853.53 L121.39 882.91 L81 881.65 L74.19 876.57 L72.11 871.41 L78.84 831.05 L123.38 815.88 L144.38 830.79 Z"
      /><path d="M144.38 830.79 L147.25 853.53 L121.39 882.91 L81 881.65 L74.19 876.57 L72.11 871.41 L78.84 831.05 L123.38 815.88 L144.38 830.79 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M356.34 208.67 L332.76 206.54 L313.79 239.76 L332.99 254.75 L360.21 248.17 L356.34 208.67 Z"
      /><path d="M356.34 208.67 L332.76 206.54 L313.79 239.76 L332.99 254.75 L360.21 248.17 L356.34 208.67 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1353.6801 457.3 L1325.74 474.37 L1343.39 515.17 L1344.66 515.81 L1380.76 501.69 L1386.13 484.95 L1353.6801 457.3 Z"
      /><path d="M1353.6801 457.3 L1325.74 474.37 L1343.39 515.17 L1344.66 515.81 L1380.76 501.69 L1386.13 484.95 L1353.6801 457.3 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M941.73 271.16 L904.99 256.18 L887.23 280.4 L899.26 303.45 L919.47 307.06 L942.13 273.59 L941.73 271.16 Z"
      /><path d="M941.73 271.16 L904.99 256.18 L887.23 280.4 L899.26 303.45 L919.47 307.06 L942.13 273.59 L941.73 271.16 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1396.64 160.23 L1376.01 127.21 L1349.73 128.01 L1343.85 166.16 L1358.66 177.07 L1396.53 160.83 L1396.64 160.23 Z"
      /><path d="M1396.64 160.23 L1376.01 127.21 L1349.73 128.01 L1343.85 166.16 L1358.66 177.07 L1396.53 160.83 L1396.64 160.23 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M139.94 402.42 L160.69 427.88 L125.38 460.08 L116.34 459.83 L100.48 419.51 L139.94 402.42 Z"
      /><path d="M139.94 402.42 L160.69 427.88 L125.38 460.08 L116.34 459.83 L100.48 419.51 L139.94 402.42 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M921.15 450.84 L910.29 455.31 L899.95 498.36 L919.3 510.83 L951.33 501.24 L960.92 475.28 L921.15 450.84 Z"
      /><path d="M921.15 450.84 L910.29 455.31 L899.95 498.36 L919.3 510.83 L951.33 501.24 L960.92 475.28 L921.15 450.84 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M1488.02 1020.63 L1455.34 1052.53 L1456.4 1080 L1520.3 1080 L1520.9301 1038.36 L1488.02 1020.63 Z"
      /><path d="M1488.02 1020.63 L1455.34 1052.53 L1456.4 1080 L1520.3 1080 L1520.9301 1038.36 L1488.02 1020.63 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1901.87 49.45 L1879.78 73.59 L1883.78 92.87 L1920 102 L1920 50.2 L1901.87 49.45 Z"
      /><path d="M1901.87 49.45 L1879.78 73.59 L1883.78 92.87 L1920 102 L1920 50.2 L1901.87 49.45 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1111.26 219.53 L1125.11 246.75 L1118.59 263.76 L1089.85 272.08 L1068.66 249.97 L1075.67 228.14 L1111.26 219.53 Z"
      /><path d="M1111.26 219.53 L1125.11 246.75 L1118.59 263.76 L1089.85 272.08 L1068.66 249.97 L1075.67 228.14 L1111.26 219.53 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1552.8 836.35 L1583.47 868.37 L1581.84 873.78 L1548.49 890.21 L1530.03 879.33 L1530.29 843.66 L1552.8 836.35 Z"
      /><path d="M1552.8 836.35 L1583.47 868.37 L1581.84 873.78 L1548.49 890.21 L1530.03 879.33 L1530.29 843.66 L1552.8 836.35 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1179.03 87.59 L1180.89 91.62 L1164.64 124.03 L1134.52 122.63 L1125.02 103.95 L1149.1801 78.26 L1179.03 87.59 Z"
      /><path d="M1179.03 87.59 L1180.89 91.62 L1164.64 124.03 L1134.52 122.63 L1125.02 103.95 L1149.1801 78.26 L1179.03 87.59 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M185.91 293.31 L213.77 315.16 L208.74 341.01 L185.14 350.2 L160.07 327.09 L164.2 303.86 L185.91 293.31 Z"
      /><path d="M185.91 293.31 L213.77 315.16 L208.74 341.01 L185.14 350.2 L160.07 327.09 L164.2 303.86 L185.91 293.31 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 975.4 L1876.58 972.05 L1875.39 1007.75 L1920 1015.5 L1920 975.4 Z"
      /><path d="M1920 975.4 L1876.58 972.05 L1875.39 1007.75 L1920 1015.5 L1920 975.4 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M872.35 939.1 L914.2 944.68 L915.26 970.5 L878.6 993.78 L872.5 990.99 L860.07 961.8 L872.35 939.1 Z"
      /><path d="M872.35 939.1 L914.2 944.68 L915.26 970.5 L878.6 993.78 L872.5 990.99 L860.07 961.8 L872.35 939.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1639.16 379.22 L1630.79 391.64 L1587.75 393.02 L1576.59 378.5 L1585.96 348.11 L1619 339.09 L1639.16 379.22 Z"
      /><path d="M1639.16 379.22 L1630.79 391.64 L1587.75 393.02 L1576.59 378.5 L1585.96 348.11 L1619 339.09 L1639.16 379.22 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1713.1 765.22 L1676 762.72 L1664.47 776.24 L1664.6899 792.94 L1694.37 815.1 L1712.6 808.1 L1713.1 765.22 Z"
      /><path d="M1713.1 765.22 L1676 762.72 L1664.47 776.24 L1664.6899 792.94 L1694.37 815.1 L1712.6 808.1 L1713.1 765.22 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M919.85 546.25 L949.33 557.48 L955.04 577.23 L938.43 597.59 L906.46 596.44 L899.01 560.14 L919.85 546.25 Z"
      /><path d="M919.85 546.25 L949.33 557.48 L955.04 577.23 L938.43 597.59 L906.46 596.44 L899.01 560.14 L919.85 546.25 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M1884.73 700.3 L1867.6 670.91 L1833.6801 681.29 L1826.96 701.99 L1862.46 728.25 L1868.66 727.1 L1884.73 700.3 Z"
      /><path d="M1884.73 700.3 L1867.6 670.91 L1833.6801 681.29 L1826.96 701.99 L1862.46 728.25 L1868.66 727.1 L1884.73 700.3 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1236.1801 961.05 L1218.05 972.94 L1214.66 995.02 L1247.41 1018.45 L1258.26 1013.71 L1267.83 975.62 L1236.1801 961.05 Z"
      /><path d="M1236.1801 961.05 L1218.05 972.94 L1214.66 995.02 L1247.41 1018.45 L1258.26 1013.71 L1267.83 975.62 L1236.1801 961.05 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1183.08 194.23 L1167.9 164.4 L1137.1801 168.66 L1127.17 196.34 L1170.8 215.28 L1183.08 194.23 Z"
      /><path d="M1183.08 194.23 L1167.9 164.4 L1137.1801 168.66 L1127.17 196.34 L1170.8 215.28 L1183.08 194.23 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M332.76 206.54 L316.01 187.35 L288.99 201.16 L288.56 228.92 L302.9 240.59 L313.79 239.76 L332.76 206.54 Z"
      /><path d="M332.76 206.54 L316.01 187.35 L288.99 201.16 L288.56 228.92 L302.9 240.59 L313.79 239.76 L332.76 206.54 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1291.36 1029.33 L1258.26 1013.71 L1247.41 1018.45 L1239.04 1036.76 L1264.6 1080 L1277.4 1080 L1291.36 1029.33 Z"
      /><path d="M1291.36 1029.33 L1258.26 1013.71 L1247.41 1018.45 L1239.04 1036.76 L1264.6 1080 L1277.4 1080 L1291.36 1029.33 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1234.0601 58.59 L1235.92 76 L1203.64 100.69 L1180.89 91.62 L1179.03 87.59 L1188.74 62.03 L1234.0601 58.59 Z"
      /><path d="M1234.0601 58.59 L1235.92 76 L1203.64 100.69 L1180.89 91.62 L1179.03 87.59 L1188.74 62.03 L1234.0601 58.59 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M979.53 429.52 L969.66 418.72 L933.12 420.38 L921.15 450.84 L960.92 475.28 L966.19 472.72 L979.53 429.52 Z"
      /><path d="M979.53 429.52 L969.66 418.72 L933.12 420.38 L921.15 450.84 L960.92 475.28 L966.19 472.72 L979.53 429.52 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M1308.4399 878.52 L1280.14 867.75 L1257.53 882.86 L1262.11 918.05 L1285.3101 928.5 L1300.1801 922.31 L1308.4399 878.52 Z"
      /><path d="M1308.4399 878.52 L1280.14 867.75 L1257.53 882.86 L1262.11 918.05 L1285.3101 928.5 L1300.1801 922.31 L1308.4399 878.52 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M931.61 843.01 L945.38 879.16 L914.58 897.03 L897.3 889.54 L894.98 844.17 L900.52 839.99 L931.61 843.01 Z"
      /><path d="M931.61 843.01 L945.38 879.16 L914.58 897.03 L897.3 889.54 L894.98 844.17 L900.52 839.99 L931.61 843.01 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1672.39 896.15 L1686.6801 923.82 L1655.11 957.31 L1641.1899 955.33 L1625.61 910.04 L1643.37 891.75 L1672.39 896.15 Z"
      /><path d="M1672.39 896.15 L1686.6801 923.82 L1655.11 957.31 L1641.1899 955.33 L1625.61 910.04 L1643.37 891.75 L1672.39 896.15 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M489.98 985.88 L511.02 987.63 L524.32 1007.81 L519.06 1032.0601 L481.43 1037.61 L463.98 1020.59 L489.98 985.88 Z"
      /><path d="M489.98 985.88 L511.02 987.63 L524.32 1007.81 L519.06 1032.0601 L481.43 1037.61 L463.98 1020.59 L489.98 985.88 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 930.4 L1920 975.4 L1876.58 972.05 L1875.54 970.71 L1889.8199 930.15 L1920 930.4 Z"
      /><path d="M1920 930.4 L1920 975.4 L1876.58 972.05 L1875.54 970.71 L1889.8199 930.15 L1920 930.4 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1270.35 783.27 L1230.4 791.58 L1227.92 828.96 L1230.13 831.05 L1274.58 833.23 L1289.9 814.35 L1270.35 783.27 Z"
      /><path d="M1270.35 783.27 L1230.4 791.58 L1227.92 828.96 L1230.13 831.05 L1274.58 833.23 L1289.9 814.35 L1270.35 783.27 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M81.71 62.36 L50.45 77.12 L70.44 112.18 L76.99 112.21 L102.48 88.92 L81.71 62.36 Z"
      /><path d="M81.71 62.36 L50.45 77.12 L70.44 112.18 L76.99 112.21 L102.48 88.92 L81.71 62.36 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1853 391.78 L1869.71 405.13 L1862.89 430.23 L1828.1801 440.17 L1810.09 425.14 L1809.42 397.88 L1811.33 396.03 L1853 391.78 Z"
      /><path d="M1853 391.78 L1869.71 405.13 L1862.89 430.23 L1828.1801 440.17 L1810.09 425.14 L1809.42 397.88 L1811.33 396.03 L1853 391.78 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M998.67 805.52 L976.48 776.41 L958.56 776.81 L941.32 796.47 L948.88 824.39 L980.08 830.88 L998.67 805.52 Z"
      /><path d="M998.67 805.52 L976.48 776.41 L958.56 776.81 L941.32 796.47 L948.88 824.39 L980.08 830.88 L998.67 805.52 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1920 362 L1920 304.9 L1889.04 306.35 L1878.16 346.08 L1898.47 362.06 L1920 362 Z"
      /><path d="M1920 362 L1920 304.9 L1889.04 306.35 L1878.16 346.08 L1898.47 362.06 L1920 362 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1804.05 508.7 L1769.09 511.96 L1758.04 536.89 L1760.2 541.89 L1797.5601 554.74 L1818.03 537.28 L1804.05 508.7 Z"
      /><path d="M1804.05 508.7 L1769.09 511.96 L1758.04 536.89 L1760.2 541.89 L1797.5601 554.74 L1818.03 537.28 L1804.05 508.7 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M301.57 327.21 L263.24 316.12 L251.75 355.45 L276.11 373.27 L285.58 371.81 L305.67 336.38 L301.57 327.21 Z"
      /><path d="M301.57 327.21 L263.24 316.12 L251.75 355.45 L276.11 373.27 L285.58 371.81 L305.67 336.38 L301.57 327.21 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1165.22 1045.87 L1153.55 1038.74 L1119.85 1053.75 L1120.4 1080 L1168.3 1080 L1165.22 1045.87 Z"
      /><path d="M1165.22 1045.87 L1153.55 1038.74 L1119.85 1053.75 L1120.4 1080 L1168.3 1080 L1165.22 1045.87 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M514.29 851.73 L523.02 855.61 L538.17 883.31 L529.74 907.42 L512.72 915.98 L485.5 893.6 L499.31 857.31 L514.29 851.73 Z"
      /><path d="M514.29 851.73 L523.02 855.61 L538.17 883.31 L529.74 907.42 L512.72 915.98 L485.5 893.6 L499.31 857.31 L514.29 851.73 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M337.43 869.88 L314.73 906.87 L297.27 905.55 L275.64 869.04 L280.97 856.45 L314.76 849.93 L337.43 869.88 Z"
      /><path d="M337.43 869.88 L314.73 906.87 L297.27 905.55 L275.64 869.04 L280.97 856.45 L314.76 849.93 L337.43 869.88 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M326.25 951.16 L359.87 974.15 L359.82 987.3 L338.31 1008.3 L301.79 990.77 L302.93 965.68 L326.25 951.16 Z"
      /><path d="M326.25 951.16 L359.87 974.15 L359.82 987.3 L338.31 1008.3 L301.79 990.77 L302.93 965.68 L326.25 951.16 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1578.02 583.8 L1551.83 616.65 L1577.55 635.02 L1598.5 628.74 L1606.12 599.03 L1578.02 583.8 Z"
      /><path d="M1578.02 583.8 L1551.83 616.65 L1577.55 635.02 L1598.5 628.74 L1606.12 599.03 L1578.02 583.8 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M681.1 471.06 L668.51 463.4 L639.61 476.76 L650.16 522.05 L686.54 509.02 L681.1 471.06 Z"
      /><path d="M681.1 471.06 L668.51 463.4 L639.61 476.76 L650.16 522.05 L686.54 509.02 L681.1 471.06 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M499.24 166.04 L523.42 187.06 L522.29 218.74 L512.13 230.52 L471.26 216.3 L470.27 187.93 L499.24 166.04 Z"
      /><path d="M499.24 166.04 L523.42 187.06 L522.29 218.74 L512.13 230.52 L471.26 216.3 L470.27 187.93 L499.24 166.04 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1531.12 332.34 L1509.9 306.75 L1488.3101 307.47 L1465.2 341.71 L1482.1899 366.03 L1524.1899 355.32 L1531.12 332.34 Z"
      /><path d="M1531.12 332.34 L1509.9 306.75 L1488.3101 307.47 L1465.2 341.71 L1482.1899 366.03 L1524.1899 355.32 L1531.12 332.34 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M125.38 460.08 L116.34 459.83 L99.28 476.33 L108.6 517.2 L129.38 523.35 L164.76 495.83 L165.34 493.73 L125.38 460.08 Z"
      /><path d="M125.38 460.08 L116.34 459.83 L99.28 476.33 L108.6 517.2 L129.38 523.35 L164.76 495.83 L165.34 493.73 L125.38 460.08 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 488.6 L1891.08 491.03 L1880.33 511.17 L1895.4301 535.28 L1920 535.8 L1920 488.6 Z"
      /><path d="M1920 488.6 L1891.08 491.03 L1880.33 511.17 L1895.4301 535.28 L1920 535.8 L1920 488.6 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M489.98 985.88 L469.09 955.65 L432.78 984.26 L457.29 1019.99 L463.98 1020.59 L489.98 985.88 Z"
      /><path d="M489.98 985.88 L469.09 955.65 L432.78 984.26 L457.29 1019.99 L463.98 1020.59 L489.98 985.88 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M527.33 1043 L565.94 1043 L572.9 1080 L523.1 1080 L527.33 1043 Z"
      /><path d="M527.33 1043 L565.94 1043 L572.9 1080 L523.1 1080 L527.33 1043 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1126.53 579.04 L1110.45 612.58 L1125.02 634.37 L1147.48 636.09 L1166.3 613.19 L1151.22 582 L1126.53 579.04 Z"
      /><path d="M1126.53 579.04 L1110.45 612.58 L1125.02 634.37 L1147.48 636.09 L1166.3 613.19 L1151.22 582 L1126.53 579.04 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M415.2 498.51 L379.93 504.84 L371.18 519.93 L397.2 546.84 L435.72 531.43 L415.2 498.51 Z"
      /><path d="M415.2 498.51 L379.93 504.84 L371.18 519.93 L397.2 546.84 L435.72 531.43 L415.2 498.51 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 753.5 L1920 698.2 L1884.73 700.3 L1868.66 727.1 L1898.05 754.18 L1920 753.5 Z"
      /><path d="M1920 753.5 L1920 698.2 L1884.73 700.3 L1868.66 727.1 L1898.05 754.18 L1920 753.5 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1100.0601 894.58 L1075.4301 927.39 L1091.21 945.14 L1133.1899 934.15 L1133.7 932.8 L1119.51 898.27 L1100.0601 894.58 Z"
      /><path d="M1100.0601 894.58 L1075.4301 927.39 L1091.21 945.14 L1133.1899 934.15 L1133.7 932.8 L1119.51 898.27 L1100.0601 894.58 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M864.87 842.26 L845.67 865.35 L870.53 899.39 L897.3 889.54 L894.98 844.17 L864.87 842.26 Z"
      /><path d="M864.87 842.26 L845.67 865.35 L870.53 899.39 L897.3 889.54 L894.98 844.17 L864.87 842.26 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M61.75 776.75 L42.15 762.81 L0 769.8 L0 825.7 L59.63 808.74 L61.75 776.75 Z"
      /><path d="M61.75 776.75 L42.15 762.81 L0 769.8 L0 825.7 L59.63 808.74 L61.75 776.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1442.35 338.01 L1432.45 289.08 L1397.41 293.45 L1386.1801 326.64 L1424.74 348.3 L1442.35 338.01 Z"
      /><path d="M1442.35 338.01 L1432.45 289.08 L1397.41 293.45 L1386.1801 326.64 L1424.74 348.3 L1442.35 338.01 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1665.4 187.98 L1677.91 193.05 L1682.29 236.85 L1654.2 246.08 L1641.37 235.61 L1645.08 198.8 L1665.4 187.98 Z"
      /><path d="M1665.4 187.98 L1677.91 193.05 L1682.29 236.85 L1654.2 246.08 L1641.37 235.61 L1645.08 198.8 L1665.4 187.98 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1066.3 774.35 L1032.83 779.36 L1019.72 803.99 L1038.8 827.94 L1076.67 818.33 L1082.64 804.75 L1066.3 774.35 Z"
      /><path d="M1066.3 774.35 L1032.83 779.36 L1019.72 803.99 L1038.8 827.94 L1076.67 818.33 L1082.64 804.75 L1066.3 774.35 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M560.34 838.95 L579.39 862.48 L574.09 878.67 L538.17 883.31 L523.02 855.61 L560.34 838.95 Z"
      /><path d="M560.34 838.95 L579.39 862.48 L574.09 878.67 L538.17 883.31 L523.02 855.61 L560.34 838.95 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1401.33 908.48 L1432.03 909.61 L1435.6899 954.1 L1430.4399 959.72 L1387.1 951.67 L1382.79 941.89 L1401.33 908.48 Z"
      /><path d="M1401.33 908.48 L1432.03 909.61 L1435.6899 954.1 L1430.4399 959.72 L1387.1 951.67 L1382.79 941.89 L1401.33 908.48 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M434.33 670.95 L427.02 701.99 L401.54 708.16 L377.17 681.08 L384.14 662.38 L414.83 652.42 L434.33 670.95 Z"
      /><path d="M434.33 670.95 L427.02 701.99 L401.54 708.16 L377.17 681.08 L384.14 662.38 L414.83 652.42 L434.33 670.95 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M308.05 751.12 L316.62 760.06 L305.36 797.85 L284.77 801.54 L253.71 770.18 L255.54 760.6 L262.14 753.6 L308.05 751.12 Z"
      /><path d="M308.05 751.12 L316.62 760.06 L305.36 797.85 L284.77 801.54 L253.71 770.18 L255.54 760.6 L262.14 753.6 L308.05 751.12 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M275.98 132.95 L279.8 154.9 L262.87 177.8 L226.08 164.11 L225.9 163.84 L252.83 121.47 L275.98 132.95 Z"
      /><path d="M275.98 132.95 L279.8 154.9 L262.87 177.8 L226.08 164.11 L225.9 163.84 L252.83 121.47 L275.98 132.95 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M209.08 220.61 L175.47 250.2 L191.06 273.87 L227.75 263.29 L209.08 220.61 Z"
      /><path d="M209.08 220.61 L175.47 250.2 L191.06 273.87 L227.75 263.29 L209.08 220.61 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1063.17 84.42 L1091.0601 103.39 L1081.42 130.1 L1044.47 128.92 L1041.99 101.03 L1063.17 84.42 Z"
      /><path d="M1063.17 84.42 L1091.0601 103.39 L1081.42 130.1 L1044.47 128.92 L1041.99 101.03 L1063.17 84.42 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1049.49 339.47 L1020.75 343.39 L1013.3 380.96 L1023.33 392.45 L1054.03 393.2 L1064.1 352.9 L1049.49 339.47 Z"
      /><path d="M1049.49 339.47 L1020.75 343.39 L1013.3 380.96 L1023.33 392.45 L1054.03 393.2 L1064.1 352.9 L1049.49 339.47 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M473.44 48.47 L458.44 25.86 L418.43 38.21 L415.19 47.05 L434.71 69.75 L466.61 62.62 L473.44 48.47 Z"
      /><path d="M473.44 48.47 L458.44 25.86 L418.43 38.21 L415.19 47.05 L434.71 69.75 L466.61 62.62 L473.44 48.47 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1186.78 954.04 L1218.05 972.94 L1214.66 995.02 L1194.54 1007.32 L1170.48 994.51 L1168.08 968.97 L1186.78 954.04 Z"
      /><path d="M1186.78 954.04 L1218.05 972.94 L1214.66 995.02 L1194.54 1007.32 L1170.48 994.51 L1168.08 968.97 L1186.78 954.04 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M982.07 334.86 L966.56 319.17 L933.34 328.14 L929.17 343.39 L947.36 369.3 L968.88 372.04 L982.07 334.86 Z"
      /><path d="M982.07 334.86 L966.56 319.17 L933.34 328.14 L929.17 343.39 L947.36 369.3 L968.88 372.04 L982.07 334.86 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M262.87 177.8 L226.08 164.11 L218.3 211.75 L245.91 214.63 L265.5 187.6 L262.87 177.8 Z"
      /><path d="M262.87 177.8 L226.08 164.11 L218.3 211.75 L245.91 214.63 L265.5 187.6 L262.87 177.8 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M676.72 978.29 L708.99 987.94 L703.79 1028.97 L692.2 1035.17 L665.55 1028.35 L657.94 1003.58 L676.72 978.29 Z"
      /><path d="M676.72 978.29 L708.99 987.94 L703.79 1028.97 L692.2 1035.17 L665.55 1028.35 L657.94 1003.58 L676.72 978.29 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1619.58 968.91 L1580.3 948.58 L1552.85 991.24 L1557.6 1005.65 L1612.27 1003.45 L1619.58 968.91 Z"
      /><path d="M1619.58 968.91 L1580.3 948.58 L1552.85 991.24 L1557.6 1005.65 L1612.27 1003.45 L1619.58 968.91 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M147.25 853.53 L121.39 882.91 L145.41 926.94 L183.95 902.17 L183.41 873.91 L147.25 853.53 Z"
      /><path d="M147.25 853.53 L121.39 882.91 L145.41 926.94 L183.95 902.17 L183.41 873.91 L147.25 853.53 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M90.71 414.15 L63.02 421.69 L52.48 449.94 L62.68 473.18 L99.28 476.33 L116.34 459.83 L100.48 419.51 L90.71 414.15 Z"
      /><path d="M90.71 414.15 L63.02 421.69 L52.48 449.94 L62.68 473.18 L99.28 476.33 L116.34 459.83 L100.48 419.51 L90.71 414.15 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M441.53 533.45 L435.72 531.43 L397.2 546.84 L393.92 579.01 L438.25 579.34 L446.53 541.53 L441.53 533.45 Z"
      /><path d="M441.53 533.45 L435.72 531.43 L397.2 546.84 L393.92 579.01 L438.25 579.34 L446.53 541.53 L441.53 533.45 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1401.33 908.48 L1382.79 941.89 L1347.55 928.47 L1351.87 893.48 L1383.88 882.02 L1401.33 908.48 Z"
      /><path d="M1401.33 908.48 L1382.79 941.89 L1347.55 928.47 L1351.87 893.48 L1383.88 882.02 L1401.33 908.48 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1599.71 40.65 L1584.79 54.22 L1584.61 79.64 L1630.3101 95.66 L1646.73 59.3 L1640.55 49.3 L1599.71 40.65 Z"
      /><path d="M1599.71 40.65 L1584.79 54.22 L1584.61 79.64 L1630.3101 95.66 L1646.73 59.3 L1640.55 49.3 L1599.71 40.65 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M0 710.2 L43.64 714.75 L42.15 762.81 L0 769.8 L0 710.2 Z"
      /><path d="M0 710.2 L43.64 714.75 L42.15 762.81 L0 769.8 L0 710.2 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M448.01 312.51 L425.28 339.7 L442.59 373.1 L442.7 373.13 L469.9 360.81 L479.87 334.79 L448.01 312.51 Z"
      /><path d="M448.01 312.51 L425.28 339.7 L442.59 373.1 L442.7 373.13 L469.9 360.81 L479.87 334.79 L448.01 312.51 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1601.5 854.96 L1634.14 861.21 L1643.37 891.75 L1625.61 910.04 L1601.11 908.48 L1581.84 873.78 L1583.47 868.37 L1601.5 854.96 Z"
      /><path d="M1601.5 854.96 L1634.14 861.21 L1643.37 891.75 L1625.61 910.04 L1601.11 908.48 L1581.84 873.78 L1583.47 868.37 L1601.5 854.96 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1895.4301 535.28 L1879.51 554.77 L1884.54 576.37 L1920 582.5 L1920 535.8 L1895.4301 535.28 Z"
      /><path d="M1895.4301 535.28 L1879.51 554.77 L1884.54 576.37 L1920 582.5 L1920 535.8 L1895.4301 535.28 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M56.14 252.55 L79.67 283.25 L64.57 301.08 L36.19 290.19 L30.71 271.2 L44.7 253.81 L56.14 252.55 Z"
      /><path d="M56.14 252.55 L79.67 283.25 L64.57 301.08 L36.19 290.19 L30.71 271.2 L44.7 253.81 L56.14 252.55 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M248.47 113.3 L252.83 121.47 L225.9 163.84 L207.23 156.78 L196.81 135.13 L209.93 112.07 L248.47 113.3 Z"
      /><path d="M248.47 113.3 L252.83 121.47 L225.9 163.84 L207.23 156.78 L196.81 135.13 L209.93 112.07 L248.47 113.3 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M368.56 52.99 L385.55 58.8 L397.34 106.07 L383.97 117.24 L364.01 116.12 L342.59 90.3 L352.34 59.64 L368.56 52.99 Z"
      /><path d="M368.56 52.99 L385.55 58.8 L397.34 106.07 L383.97 117.24 L364.01 116.12 L342.59 90.3 L352.34 59.64 L368.56 52.99 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1392.92 858.01 L1391.61 858.61 L1383.88 882.02 L1401.33 908.48 L1432.03 909.61 L1445.15 898.22 L1446.63 892.37 L1437.03 869.46 L1392.92 858.01 Z"
      /><path d="M1392.92 858.01 L1391.61 858.61 L1383.88 882.02 L1401.33 908.48 L1432.03 909.61 L1445.15 898.22 L1446.63 892.37 L1437.03 869.46 L1392.92 858.01 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M101.48 710.87 L143.18 728.36 L145.37 759.14 L120.99 777.28 L89.28 763.43 L91.58 717.52 L101.48 710.87 Z"
      /><path d="M101.48 710.87 L143.18 728.36 L145.37 759.14 L120.99 777.28 L89.28 763.43 L91.58 717.52 L101.48 710.87 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M451.17 250.84 L474.37 275.04 L447.68 310.39 L418.45 287.56 L421.8 265.31 L451.17 250.84 Z"
      /><path d="M451.17 250.84 L474.37 275.04 L447.68 310.39 L418.45 287.56 L421.8 265.31 L451.17 250.84 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M342.02 562.92 L347.82 574.24 L330.37 608.73 L290.51 600.39 L286.91 590.23 L306.5 552.95 L342.02 562.92 Z"
      /><path d="M342.02 562.92 L347.82 574.24 L330.37 608.73 L290.51 600.39 L286.91 590.23 L306.5 552.95 L342.02 562.92 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M582.98 305.27 L549.22 275.88 L526.15 301.36 L543.75 336.54 L551.09 337.73 L582.98 305.27 Z"
      /><path d="M582.98 305.27 L549.22 275.88 L526.15 301.36 L543.75 336.54 L551.09 337.73 L582.98 305.27 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1424.98 241.12 L1403.2 235.67 L1378.1801 270.19 L1397.41 293.45 L1432.45 289.08 L1437.24 283.59 L1424.98 241.12 Z"
      /><path d="M1424.98 241.12 L1403.2 235.67 L1378.1801 270.19 L1397.41 293.45 L1432.45 289.08 L1437.24 283.59 L1424.98 241.12 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M32.9 0 L0 0 L0 46.1 L33.21 44.77 L39.5 36.03 L32.9 0 Z"
      /><path d="M32.9 0 L0 0 L0 46.1 L33.21 44.77 L39.5 36.03 L32.9 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1858.49 144.87 L1883.54 184.29 L1871.84 207.17 L1859.64 212.79 L1843.1801 208.4 L1825.73 176.97 L1858.49 144.87 Z"
      /><path d="M1858.49 144.87 L1883.54 184.29 L1871.84 207.17 L1859.64 212.79 L1843.1801 208.4 L1825.73 176.97 L1858.49 144.87 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1895.4301 535.28 L1880.33 511.17 L1854.88 513.74 L1839.72 541.25 L1841.55 543.97 L1879.51 554.77 L1895.4301 535.28 Z"
      /><path d="M1895.4301 535.28 L1880.33 511.17 L1854.88 513.74 L1839.72 541.25 L1841.55 543.97 L1879.51 554.77 L1895.4301 535.28 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M995.1 0 L1054.4 0 L1035.88 37.08 L1000.83 28.15 L995.1 0 Z"
      /><path d="M995.1 0 L1054.4 0 L1035.88 37.08 L1000.83 28.15 L995.1 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M231.31 264.78 L234.78 304.04 L213.77 315.16 L185.91 293.31 L191.06 273.87 L227.75 263.29 L231.31 264.78 Z"
      /><path d="M231.31 264.78 L234.78 304.04 L213.77 315.16 L185.91 293.31 L191.06 273.87 L227.75 263.29 L231.31 264.78 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1086.6 406.73 L1066.8199 406.2 L1049.77 448.68 L1063.16 463.82 L1103.6899 456.55 L1111.52 433.34 L1086.6 406.73 Z"
      /><path d="M1086.6 406.73 L1066.8199 406.2 L1049.77 448.68 L1063.16 463.82 L1103.6899 456.55 L1111.52 433.34 L1086.6 406.73 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1495.33 614.46 L1488.85 612.37 L1464.5601 645.32 L1469.23 661.89 L1496.15 670.39 L1516.9 656.49 L1495.33 614.46 Z"
      /><path d="M1495.33 614.46 L1488.85 612.37 L1464.5601 645.32 L1469.23 661.89 L1496.15 670.39 L1516.9 656.49 L1495.33 614.46 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M77 0 L116.8 0 L114.54 37.01 L84.8 46.12 L73.08 32.67 L77 0 Z"
      /><path d="M77 0 L116.8 0 L114.54 37.01 L84.8 46.12 L73.08 32.67 L77 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1040.0699 291.49 L1056.8 304.97 L1049.49 339.47 L1020.75 343.39 L1008.16 332.35 L1014.29 297.03 L1040.0699 291.49 Z"
      /><path d="M1040.0699 291.49 L1056.8 304.97 L1049.49 339.47 L1020.75 343.39 L1008.16 332.35 L1014.29 297.03 L1040.0699 291.49 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M991.33 612.93 L1022.44 621.49 L1028.23 645.64 L993.99 670.18 L971.75 633.14 L991.33 612.93 Z"
      /><path d="M991.33 612.93 L1022.44 621.49 L1028.23 645.64 L993.99 670.18 L971.75 633.14 L991.33 612.93 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1700.05 648.99 L1679.0699 648.03 L1668.29 660.2 L1674.28 687.65 L1694.49 696.82 L1715.08 669.86 L1700.05 648.99 Z"
      /><path d="M1700.05 648.99 L1679.0699 648.03 L1668.29 660.2 L1674.28 687.65 L1694.49 696.82 L1715.08 669.86 L1700.05 648.99 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M467.78 897.01 L453.37 930.28 L425.63 928.74 L414.21 913.51 L418.35 886.73 L443.67 875.98 L467.78 897.01 Z"
      /><path d="M467.78 897.01 L453.37 930.28 L425.63 928.74 L414.21 913.51 L418.35 886.73 L443.67 875.98 L467.78 897.01 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M669.86 606.61 L639.38 583.65 L629.74 586.07 L616.99 622.23 L640.93 644.84 L661.97 640.38 L669.86 606.61 Z"
      /><path d="M669.86 606.61 L639.38 583.65 L629.74 586.07 L616.99 622.23 L640.93 644.84 L661.97 640.38 L669.86 606.61 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M717.95 983.19 L752.37 1001.03 L753.92 1025.98 L730.61 1039.0601 L703.79 1028.97 L708.99 987.94 L717.95 983.19 Z"
      /><path d="M717.95 983.19 L752.37 1001.03 L753.92 1025.98 L730.61 1039.0601 L703.79 1028.97 L708.99 987.94 L717.95 983.19 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M815.87 138.01 L795.5 129.14 L771.29 159.63 L782.12 175.02 L820.51 165.31 L815.87 138.01 Z"
      /><path d="M815.87 138.01 L795.5 129.14 L771.29 159.63 L782.12 175.02 L820.51 165.31 L815.87 138.01 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1211.77 1047.34 L1193.4 1033.36 L1165.22 1045.87 L1168.3 1080 L1209 1080 L1211.77 1047.34 Z"
      /><path d="M1211.77 1047.34 L1193.4 1033.36 L1165.22 1045.87 L1168.3 1080 L1209 1080 L1211.77 1047.34 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1269.7 324.31 L1250.73 314.49 L1223.54 331.81 L1222.4399 364.42 L1246.5601 381.9 L1256.78 379.3 L1276.92 352.59 L1269.7 324.31 Z"
      /><path d="M1269.7 324.31 L1250.73 314.49 L1223.54 331.81 L1222.4399 364.42 L1246.5601 381.9 L1256.78 379.3 L1276.92 352.59 L1269.7 324.31 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M48.21 496.29 L0 495.6 L0 546.2 L37.91 550.47 L60.04 531.31 L48.21 496.29 Z"
      /><path d="M48.21 496.29 L0 495.6 L0 546.2 L37.91 550.47 L60.04 531.31 L48.21 496.29 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M585.54 695.16 L604.12 726.32 L587.31 746.73 L550.55 738.73 L543.72 724.37 L563.86 696.82 L585.54 695.16 Z"
      /><path d="M585.54 695.16 L604.12 726.32 L587.31 746.73 L550.55 738.73 L543.72 724.37 L563.86 696.82 L585.54 695.16 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M699.7 0 L698.26 41.61 L681.36 52.39 L648.81 42.16 L650.7 0 L699.7 0 Z"
      /><path d="M699.7 0 L698.26 41.61 L681.36 52.39 L648.81 42.16 L650.7 0 L699.7 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1094.63 349.46 L1112.77 368.32 L1086.6 406.73 L1066.8199 406.2 L1054.03 393.2 L1064.1 352.9 L1094.63 349.46 Z"
      /><path d="M1094.63 349.46 L1112.77 368.32 L1086.6 406.73 L1066.8199 406.2 L1054.03 393.2 L1064.1 352.9 L1094.63 349.46 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M122.77 131.98 L150.72 153.18 L151.11 162.7 L130.63 181.81 L110.36 177.97 L98.03 150.45 L100.82 143.49 L122.77 131.98 Z"
      /><path d="M122.77 131.98 L150.72 153.18 L151.11 162.7 L130.63 181.81 L110.36 177.97 L98.03 150.45 L100.82 143.49 L122.77 131.98 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1623.71 761.78 L1664.47 776.24 L1664.6899 792.94 L1639.54 813.74 L1620.66 807.62 L1614.12 771.64 L1623.71 761.78 Z"
      /><path d="M1623.71 761.78 L1664.47 776.24 L1664.6899 792.94 L1639.54 813.74 L1620.66 807.62 L1614.12 771.64 L1623.71 761.78 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1289.8199 515.82 L1263.67 525.19 L1258.97 556.57 L1274.72 568.38 L1305.42 554.08 L1304.74 528.4 L1289.8199 515.82 Z"
      /><path d="M1289.8199 515.82 L1263.67 525.19 L1258.97 556.57 L1274.72 568.38 L1305.42 554.08 L1304.74 528.4 L1289.8199 515.82 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M389.85 604.2 L419.65 627.06 L414.83 652.42 L384.14 662.38 L363.82 632.41 L389.85 604.2 Z"
      /><path d="M389.85 604.2 L419.65 627.06 L414.83 652.42 L384.14 662.38 L363.82 632.41 L389.85 604.2 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1070.17 178.46 L1058.5 204.06 L1034.9301 207.71 L1013.26 177.72 L1014.77 171.79 L1035.97 154.78 L1070.17 178.46 Z"
      /><path d="M1070.17 178.46 L1058.5 204.06 L1034.9301 207.71 L1013.26 177.72 L1014.77 171.79 L1035.97 154.78 L1070.17 178.46 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1185.37 670.21 L1164.4399 669.08 L1144.88 689.96 L1147.16 714.99 L1168.15 731.16 L1196.42 721.82 L1204.77 697.74 L1185.37 670.21 Z"
      /><path d="M1185.37 670.21 L1164.4399 669.08 L1144.88 689.96 L1147.16 714.99 L1168.15 731.16 L1196.42 721.82 L1204.77 697.74 L1185.37 670.21 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M270.79 931.66 L237.46 906.55 L212.51 920.33 L210.58 951.25 L244.09 968.82 L271.25 944.86 L270.79 931.66 Z"
      /><path d="M270.79 931.66 L237.46 906.55 L212.51 920.33 L210.58 951.25 L244.09 968.82 L271.25 944.86 L270.79 931.66 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1587.55 521.9 L1553.4399 524.47 L1550.25 559.79 L1574.97 573.44 L1602.1801 542.44 L1587.55 521.9 Z"
      /><path d="M1587.55 521.9 L1553.4399 524.47 L1550.25 559.79 L1574.97 573.44 L1602.1801 542.44 L1587.55 521.9 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1257.53 882.86 L1233.39 874.91 L1213.75 886.6 L1217.38 920.1 L1236.63 931.17 L1262.11 918.05 L1257.53 882.86 Z"
      /><path d="M1257.53 882.86 L1233.39 874.91 L1213.75 886.6 L1217.38 920.1 L1236.63 931.17 L1262.11 918.05 L1257.53 882.86 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M305.36 797.85 L323.56 814.24 L314.76 849.93 L280.97 856.45 L267.97 830.51 L284.77 801.54 L305.36 797.85 Z"
      /><path d="M305.36 797.85 L323.56 814.24 L314.76 849.93 L280.97 856.45 L267.97 830.51 L284.77 801.54 L305.36 797.85 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1527.22 935.08 L1522.3 971.41 L1491.51 980.97 L1472.98 951.28 L1482.12 927.92 L1500.26 919.25 L1527.22 935.08 Z"
      /><path d="M1527.22 935.08 L1522.3 971.41 L1491.51 980.97 L1472.98 951.28 L1482.12 927.92 L1500.26 919.25 L1527.22 935.08 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1254.46 734.96 L1277.4301 760.51 L1270.35 783.27 L1230.4 791.58 L1215.47 776.05 L1221.15 747.73 L1254.46 734.96 Z"
      /><path d="M1254.46 734.96 L1277.4301 760.51 L1270.35 783.27 L1230.4 791.58 L1215.47 776.05 L1221.15 747.73 L1254.46 734.96 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1611.35 170.9 L1617.89 189.49 L1601.74 212.06 L1575.04 211.24 L1569.9 171.75 L1611.35 170.9 Z"
      /><path d="M1611.35 170.9 L1617.89 189.49 L1601.74 212.06 L1575.04 211.24 L1569.9 171.75 L1611.35 170.9 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M833.53 643.96 L857.26 653.3 L847.69 697.79 L832.16 705.26 L801.92 679.22 L804.87 660.08 L833.53 643.96 Z"
      /><path d="M833.53 643.96 L857.26 653.3 L847.69 697.79 L832.16 705.26 L801.92 679.22 L804.87 660.08 L833.53 643.96 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1168.1899 467.78 L1193.79 478.96 L1201.15 519.65 L1172.95 535.64 L1153.61 524.25 L1149.99 483.05 L1168.1899 467.78 Z"
      /><path d="M1168.1899 467.78 L1193.79 478.96 L1201.15 519.65 L1172.95 535.64 L1153.61 524.25 L1149.99 483.05 L1168.1899 467.78 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1691.84 92.85 L1739.89 104.52 L1735.51 125.18 L1704.8199 146.48 L1674.46 131.47 L1672.52 121.11 L1691.84 92.85 Z"
      /><path d="M1691.84 92.85 L1739.89 104.52 L1735.51 125.18 L1704.8199 146.48 L1674.46 131.47 L1672.52 121.11 L1691.84 92.85 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M677.35 691.73 L715.15 697.93 L724.43 726.1 L686.63 745.43 L676.55 741.08 L667.74 699.74 L677.35 691.73 Z"
      /><path d="M677.35 691.73 L715.15 697.93 L724.43 726.1 L686.63 745.43 L676.55 741.08 L667.74 699.74 L677.35 691.73 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1617.89 189.49 L1645.08 198.8 L1641.37 235.61 L1615.63 237.32 L1601.74 212.06 L1617.89 189.49 Z"
      /><path d="M1617.89 189.49 L1645.08 198.8 L1641.37 235.61 L1615.63 237.32 L1601.74 212.06 L1617.89 189.49 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M584.23 646.89 L549.13 651.42 L540.59 663.3 L563.86 696.82 L585.54 695.16 L598.66 674.42 L584.23 646.89 Z"
      /><path d="M584.23 646.89 L549.13 651.42 L540.59 663.3 L563.86 696.82 L585.54 695.16 L598.66 674.42 L584.23 646.89 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M191.45 545.43 L190.14 550.37 L142.31 558.6 L129.38 523.35 L164.76 495.83 L191.45 545.43 Z"
      /><path d="M191.45 545.43 L190.14 550.37 L142.31 558.6 L129.38 523.35 L164.76 495.83 L191.45 545.43 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M643.45 697.68 L667.74 699.74 L676.55 741.08 L644.56 755.74 L621.67 726.2 L643.45 697.68 Z"
      /><path d="M643.45 697.68 L667.74 699.74 L676.55 741.08 L644.56 755.74 L621.67 726.2 L643.45 697.68 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1602.1801 542.44 L1619.76 546.25 L1626.83 558.18 L1613.64 596.12 L1606.12 599.03 L1578.02 583.8 L1574.97 573.44 L1602.1801 542.44 Z"
      /><path d="M1602.1801 542.44 L1619.76 546.25 L1626.83 558.18 L1613.64 596.12 L1606.12 599.03 L1578.02 583.8 L1574.97 573.44 L1602.1801 542.44 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M701.55 336.31 L677.15 338.2 L658.12 375.55 L698.43 391.7 L721.04 370.37 L701.55 336.31 Z"
      /><path d="M701.55 336.31 L677.15 338.2 L658.12 375.55 L698.43 391.7 L721.04 370.37 L701.55 336.31 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M795.81 396.68 L831.79 409.55 L831.41 444.97 L811.74 455.03 L786.23 442.63 L789.71 401.09 L795.81 396.68 Z"
      /><path d="M795.81 396.68 L831.79 409.55 L831.41 444.97 L811.74 455.03 L786.23 442.63 L789.71 401.09 L795.81 396.68 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1868.66 727.1 L1862.46 728.25 L1839.4 759.4 L1857.22 787.4 L1871.04 788.85 L1898.05 754.18 L1868.66 727.1 Z"
      /><path d="M1868.66 727.1 L1862.46 728.25 L1839.4 759.4 L1857.22 787.4 L1871.04 788.85 L1898.05 754.18 L1868.66 727.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1486.61 875.81 L1503.55 889.62 L1500.26 919.25 L1482.12 927.92 L1445.15 898.22 L1446.63 892.37 L1486.61 875.81 Z"
      /><path d="M1486.61 875.81 L1503.55 889.62 L1500.26 919.25 L1482.12 927.92 L1445.15 898.22 L1446.63 892.37 L1486.61 875.81 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1889.8199 930.15 L1871.77 911.85 L1837.64 936.51 L1842.27 962.59 L1875.54 970.71 L1889.8199 930.15 Z"
      /><path d="M1889.8199 930.15 L1871.77 911.85 L1837.64 936.51 L1842.27 962.59 L1875.54 970.71 L1889.8199 930.15 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M543.72 724.37 L524.87 719.02 L494.57 738.83 L492.8 754.37 L508.48 772.43 L539.09 766.71 L550.55 738.73 L543.72 724.37 Z"
      /><path d="M543.72 724.37 L524.87 719.02 L494.57 738.83 L492.8 754.37 L508.48 772.43 L539.09 766.71 L550.55 738.73 L543.72 724.37 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M510.79 685.97 L481.39 689.46 L470.92 712.95 L494.57 738.83 L524.87 719.02 L510.79 685.97 Z"
      /><path d="M510.79 685.97 L481.39 689.46 L470.92 712.95 L494.57 738.83 L524.87 719.02 L510.79 685.97 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1353.65 708.31 L1365.7 740.73 L1359.77 751.15 L1325.1801 761.94 L1310.14 750.49 L1311.9 720.43 L1344.97 703.61 L1353.65 708.31 Z"
      /><path d="M1353.65 708.31 L1365.7 740.73 L1359.77 751.15 L1325.1801 761.94 L1310.14 750.49 L1311.9 720.43 L1344.97 703.61 L1353.65 708.31 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1647.64 702.72 L1634.17 693.12 L1611.78 695.81 L1601.1801 722.35 L1624.79 742.97 L1650.48 725.5 L1647.64 702.72 Z"
      /><path d="M1647.64 702.72 L1634.17 693.12 L1611.78 695.81 L1601.1801 722.35 L1624.79 742.97 L1650.48 725.5 L1647.64 702.72 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1245.58 480.74 L1222.38 464.89 L1193.79 478.96 L1201.15 519.65 L1213.3199 523.34 L1242.08 509.3 L1245.58 480.74 Z"
      /><path d="M1245.58 480.74 L1222.38 464.89 L1193.79 478.96 L1201.15 519.65 L1213.3199 523.34 L1242.08 509.3 L1245.58 480.74 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M589.86 140.28 L621.14 154.44 L618.34 195.17 L583.65 206.15 L561.03 171.49 L564.85 154.91 L589.86 140.28 Z"
      /><path d="M589.86 140.28 L621.14 154.44 L618.34 195.17 L583.65 206.15 L561.03 171.49 L564.85 154.91 L589.86 140.28 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M143.06 665.78 L107.18 683.97 L101.48 710.87 L143.18 728.36 L163.42 709.4 L146.23 666.74 L143.06 665.78 Z"
      /><path d="M143.06 665.78 L107.18 683.97 L101.48 710.87 L143.18 728.36 L163.42 709.4 L146.23 666.74 L143.06 665.78 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1134.52 122.63 L1122.88 147.29 L1137.1801 168.66 L1167.9 164.4 L1177.91 146.08 L1164.64 124.03 L1134.52 122.63 Z"
      /><path d="M1134.52 122.63 L1122.88 147.29 L1137.1801 168.66 L1167.9 164.4 L1177.91 146.08 L1164.64 124.03 L1134.52 122.63 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 874.1 L1920 930.4 L1889.8199 930.15 L1871.77 911.85 L1871.54 905.64 L1907.65 874.15 L1920 874.1 Z"
      /><path d="M1920 874.1 L1920 930.4 L1889.8199 930.15 L1871.77 911.85 L1871.54 905.64 L1907.65 874.15 L1920 874.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M582.98 305.27 L590.12 305.37 L612.88 329.98 L575.42 369.03 L551.09 337.73 L582.98 305.27 Z"
      /><path d="M582.98 305.27 L590.12 305.37 L612.88 329.98 L575.42 369.03 L551.09 337.73 L582.98 305.27 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1214.66 995.02 L1247.41 1018.45 L1239.04 1036.76 L1211.77 1047.34 L1193.4 1033.36 L1194.54 1007.32 L1214.66 995.02 Z"
      /><path d="M1214.66 995.02 L1247.41 1018.45 L1239.04 1036.76 L1211.77 1047.34 L1193.4 1033.36 L1194.54 1007.32 L1214.66 995.02 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M511.79 90.52 L481.54 99.1 L478.6 103.61 L479.43 132.99 L499.05 151.69 L533.77 128.71 L534.98 104.74 L511.79 90.52 Z"
      /><path d="M511.79 90.52 L481.54 99.1 L478.6 103.61 L479.43 132.99 L499.05 151.69 L533.77 128.71 L534.98 104.74 L511.79 90.52 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1141.4399 959.62 L1133.1899 934.15 L1091.21 945.14 L1090.62 969.22 L1122.3101 982.09 L1141.4399 959.62 Z"
      /><path d="M1141.4399 959.62 L1133.1899 934.15 L1091.21 945.14 L1090.62 969.22 L1122.3101 982.09 L1141.4399 959.62 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1865.0699 111.69 L1830.99 86.85 L1808.5 102.35 L1804.3199 118.91 L1858.49 144.85 L1863.37 138.52 L1865.0699 111.69 Z"
      /><path d="M1865.0699 111.69 L1830.99 86.85 L1808.5 102.35 L1804.3199 118.91 L1858.49 144.85 L1863.37 138.52 L1865.0699 111.69 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1447.8 788.39 L1471.88 812.56 L1466.95 836.74 L1450.55 841.9 L1417.76 816.16 L1447.8 788.39 Z"
      /><path d="M1447.8 788.39 L1471.88 812.56 L1466.95 836.74 L1450.55 841.9 L1417.76 816.16 L1447.8 788.39 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1598.5 628.74 L1577.55 635.02 L1571.74 667.54 L1577.45 674.82 L1596.96 677.49 L1618.72 647.15 L1598.5 628.74 Z"
      /><path d="M1598.5 628.74 L1577.55 635.02 L1571.74 667.54 L1577.45 674.82 L1596.96 677.49 L1618.72 647.15 L1598.5 628.74 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1135.65 816.87 L1129.64 844.87 L1092.49 851.62 L1076.67 818.33 L1082.64 804.75 L1119.64 796.74 L1135.65 816.87 Z"
      /><path d="M1135.65 816.87 L1129.64 844.87 L1092.49 851.62 L1076.67 818.33 L1082.64 804.75 L1119.64 796.74 L1135.65 816.87 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M260.22 632.73 L231.39 619.33 L222.48 623.62 L209.42 666.77 L239.36 680.64 L254.08 670.77 L260.22 632.73 Z"
      /><path d="M260.22 632.73 L231.39 619.33 L222.48 623.62 L209.42 666.77 L239.36 680.64 L254.08 670.77 L260.22 632.73 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M183.95 902.17 L212.51 920.33 L210.58 951.25 L188.17 965.95 L144.08 932.08 L145.41 926.94 L183.95 902.17 Z"
      /><path d="M183.95 902.17 L212.51 920.33 L210.58 951.25 L188.17 965.95 L144.08 932.08 L145.41 926.94 L183.95 902.17 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M643.45 697.68 L621.67 726.2 L604.12 726.32 L585.54 695.16 L598.66 674.42 L627.19 672.96 L643.45 697.68 Z"
      /><path d="M643.45 697.68 L621.67 726.2 L604.12 726.32 L585.54 695.16 L598.66 674.42 L627.19 672.96 L643.45 697.68 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M545.94 491.11 L530.85 475.57 L500.61 477.86 L487.61 501.21 L501.97 523.26 L523.99 523.57 L545.94 491.11 Z"
      /><path d="M545.94 491.11 L530.85 475.57 L500.61 477.86 L487.61 501.21 L501.97 523.26 L523.99 523.57 L545.94 491.11 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 0 L1920 50.2 L1901.87 49.45 L1885.8199 31.69 L1893.3 0 L1920 0 Z"
      /><path d="M1920 0 L1920 50.2 L1901.87 49.45 L1885.8199 31.69 L1893.3 0 L1920 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1359.77 751.15 L1380.71 792.56 L1363.77 805.77 L1327 792.95 L1325.1801 761.94 L1359.77 751.15 Z"
      /><path d="M1359.77 751.15 L1380.71 792.56 L1363.77 805.77 L1327 792.95 L1325.1801 761.94 L1359.77 751.15 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1100.0601 894.58 L1084.63 868.16 L1055.74 873.61 L1044.84 905.86 L1061.53 926.05 L1075.4301 927.39 L1100.0601 894.58 Z"
      /><path d="M1100.0601 894.58 L1084.63 868.16 L1055.74 873.61 L1044.84 905.86 L1061.53 926.05 L1075.4301 927.39 L1100.0601 894.58 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M851.3 0 L897.5 0 L898.41 12.65 L874.04 43.79 L861.76 43.84 L851.97 34.74 L851.3 0 Z"
      /><path d="M851.3 0 L897.5 0 L898.41 12.65 L874.04 43.79 L861.76 43.84 L851.97 34.74 L851.3 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1562.88 708.94 L1534.63 708.33 L1528.27 713.07 L1527.38 747.7 L1538.6899 757.67 L1570.73 751.87 L1579.21 727.43 L1562.88 708.94 Z"
      /><path d="M1562.88 708.94 L1534.63 708.33 L1528.27 713.07 L1527.38 747.7 L1538.6899 757.67 L1570.73 751.87 L1579.21 727.43 L1562.88 708.94 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M592.17 49.19 L603.85 93.07 L589.47 105.36 L554.16 93.59 L558.26 52.58 L592.17 49.19 Z"
      /><path d="M592.17 49.19 L603.85 93.07 L589.47 105.36 L554.16 93.59 L558.26 52.58 L592.17 49.19 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M232.17 464.38 L268.31 469.82 L274.19 494.38 L250.79 526.44 L227.9 518.33 L217.6 490.94 L232.17 464.38 Z"
      /><path d="M232.17 464.38 L268.31 469.82 L274.19 494.38 L250.79 526.44 L227.9 518.33 L217.6 490.94 L232.17 464.38 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1535.55 122.04 L1524.22 131.58 L1524.9301 148.16 L1550.15 170.6 L1566.74 168.99 L1572.36 132.14 L1535.55 122.04 Z"
      /><path d="M1535.55 122.04 L1524.22 131.58 L1524.9301 148.16 L1550.15 170.6 L1566.74 168.99 L1572.36 132.14 L1535.55 122.04 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1344.66 515.81 L1352.8101 547.97 L1322.76 566.95 L1305.42 554.08 L1304.74 528.4 L1343.39 515.17 L1344.66 515.81 Z"
      /><path d="M1344.66 515.81 L1352.8101 547.97 L1322.76 566.95 L1305.42 554.08 L1304.74 528.4 L1343.39 515.17 L1344.66 515.81 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1859.64 212.79 L1843.1801 208.4 L1814.38 231.44 L1829.28 262.87 L1860.83 255.88 L1859.64 212.79 Z"
      /><path d="M1859.64 212.79 L1843.1801 208.4 L1814.38 231.44 L1829.28 262.87 L1860.83 255.88 L1859.64 212.79 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1141.4399 959.62 L1122.3101 982.09 L1126.39 1002.39 L1147.26 1010.64 L1170.48 994.51 L1168.08 968.97 L1141.4399 959.62 Z"
      /><path d="M1141.4399 959.62 L1122.3101 982.09 L1126.39 1002.39 L1147.26 1010.64 L1170.48 994.51 L1168.08 968.97 L1141.4399 959.62 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M887.23 280.4 L861.05 276.9 L843.69 303.41 L873.73 333.95 L899.26 303.45 L887.23 280.4 Z"
      /><path d="M887.23 280.4 L861.05 276.9 L843.69 303.41 L873.73 333.95 L899.26 303.45 L887.23 280.4 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1791.29 146.19 L1759.11 159.24 L1754.21 172.13 L1765.0601 197.15 L1786.53 202.69 L1812.2 175.39 L1791.29 146.19 Z"
      /><path d="M1791.29 146.19 L1759.11 159.24 L1754.21 172.13 L1765.0601 197.15 L1786.53 202.69 L1812.2 175.39 L1791.29 146.19 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M372.4 256.04 L372.4 278.7 L342.87 298.13 L326.64 291.37 L332.99 254.75 L360.21 248.17 L372.4 256.04 Z"
      /><path d="M372.4 256.04 L372.4 278.7 L342.87 298.13 L326.64 291.37 L332.99 254.75 L360.21 248.17 L372.4 256.04 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M629.93 919.28 L627.75 918.29 L594.02 945.59 L606.17 977.75 L615.33 981.56 L645.09 952.92 L629.93 919.28 Z"
      /><path d="M629.93 919.28 L627.75 918.29 L594.02 945.59 L606.17 977.75 L615.33 981.56 L645.09 952.92 L629.93 919.28 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1433.46 760.75 L1448.1899 780.85 L1447.8 788.39 L1417.76 816.16 L1416.72 816.25 L1389.11 792.48 L1413.1801 760.19 L1433.46 760.75 Z"
      /><path d="M1433.46 760.75 L1448.1899 780.85 L1447.8 788.39 L1417.76 816.16 L1416.72 816.25 L1389.11 792.48 L1413.1801 760.19 L1433.46 760.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M642.48 212.11 L644.06 234.27 L621.86 262.32 L615.46 263.35 L579.02 240.46 L575.69 224.19 L583.65 206.15 L618.34 195.17 L642.48 212.11 Z"
      /><path d="M642.48 212.11 L644.06 234.27 L621.86 262.32 L615.46 263.35 L579.02 240.46 L575.69 224.19 L583.65 206.15 L618.34 195.17 L642.48 212.11 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1797.21 125.32 L1740.98 103.56 L1739.89 104.52 L1735.51 125.18 L1759.11 159.24 L1791.29 146.19 L1797.21 125.32 Z"
      /><path d="M1797.21 125.32 L1740.98 103.56 L1739.89 104.52 L1735.51 125.18 L1759.11 159.24 L1791.29 146.19 L1797.21 125.32 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M759.85 474.33 L789.56 498.82 L784.17 519.21 L764.23 530.54 L748.15 526.47 L732.37 495.31 L734.69 487.02 L759.85 474.33 Z"
      /><path d="M759.85 474.33 L789.56 498.82 L784.17 519.21 L764.23 530.54 L748.15 526.47 L732.37 495.31 L734.69 487.02 L759.85 474.33 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M495.46 636.55 L470.77 646.38 L463.86 663.1 L481.39 689.46 L510.79 685.97 L523.19 667.27 L495.46 636.55 Z"
      /><path d="M495.46 636.55 L470.77 646.38 L463.86 663.1 L481.39 689.46 L510.79 685.97 L523.19 667.27 L495.46 636.55 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M519.06 1032.0601 L527.33 1043 L523.1 1080 L477.8 1080 L481.43 1037.61 L519.06 1032.0601 Z"
      /><path d="M519.06 1032.0601 L527.33 1043 L523.1 1080 L477.8 1080 L481.43 1037.61 L519.06 1032.0601 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1271.65 191.72 L1253.75 172.39 L1221.03 181.57 L1216.65 188.6 L1230.9 230.56 L1242.95 231.69 L1267.59 215.7 L1271.65 191.72 Z"
      /><path d="M1271.65 191.72 L1253.75 172.39 L1221.03 181.57 L1216.65 188.6 L1230.9 230.56 L1242.95 231.69 L1267.59 215.7 L1271.65 191.72 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1613.64 596.12 L1644.1801 608.46 L1647.49 615.53 L1629.6899 647.33 L1618.72 647.15 L1598.5 628.74 L1606.12 599.03 L1613.64 596.12 Z"
      /><path d="M1613.64 596.12 L1644.1801 608.46 L1647.49 615.53 L1629.6899 647.33 L1618.72 647.15 L1598.5 628.74 L1606.12 599.03 L1613.64 596.12 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M364.81 789.89 L346.66 757.94 L316.62 760.06 L305.36 797.85 L323.56 814.24 L354.92 810.43 L364.81 789.89 Z"
      /><path d="M364.81 789.89 L346.66 757.94 L316.62 760.06 L305.36 797.85 L323.56 814.24 L354.92 810.43 L364.81 789.89 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M394.2 157.52 L430.66 165.82 L431.39 167.69 L416.65 209.85 L405.09 215.07 L371.14 197.3 L372.08 175.33 L394.2 157.52 Z"
      /><path d="M394.2 157.52 L430.66 165.82 L431.39 167.69 L416.65 209.85 L405.09 215.07 L371.14 197.3 L372.08 175.33 L394.2 157.52 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1445.15 898.22 L1432.03 909.61 L1435.6899 954.1 L1472.98 951.28 L1482.12 927.92 L1445.15 898.22 Z"
      /><path d="M1445.15 898.22 L1432.03 909.61 L1435.6899 954.1 L1472.98 951.28 L1482.12 927.92 L1445.15 898.22 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M658.12 375.55 L698.43 391.7 L700.52 417.35 L666.46 433.01 L649.22 420.63 L654.49 377.03 L658.12 375.55 Z"
      /><path d="M658.12 375.55 L698.43 391.7 L700.52 417.35 L666.46 433.01 L649.22 420.63 L654.49 377.03 L658.12 375.55 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M335.35 463.79 L370.85 468.92 L379.93 504.84 L371.18 519.93 L362.19 522.77 L322.11 502.54 L328.89 469.16 L335.35 463.79 Z"
      /><path d="M335.35 463.79 L370.85 468.92 L379.93 504.84 L371.18 519.93 L362.19 522.77 L322.11 502.54 L328.89 469.16 L335.35 463.79 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M636.76 371.08 L601.49 390.81 L603.61 419.04 L619.77 429.11 L649.22 420.63 L654.49 377.03 L636.76 371.08 Z"
      /><path d="M636.76 371.08 L601.49 390.81 L603.61 419.04 L619.77 429.11 L649.22 420.63 L654.49 377.03 L636.76 371.08 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1001.66 1012.65 L1020.45 1013.34 L1036.8101 1031.1899 L1016.5 1080 L1005 1080 L982.75 1030.75 L1001.66 1012.65 Z"
      /><path d="M1001.66 1012.65 L1020.45 1013.34 L1036.8101 1031.1899 L1016.5 1080 L1005 1080 L982.75 1030.75 L1001.66 1012.65 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M921.31 1041.76 L948.85 1052.3199 L952 1080 L900.1 1080 L900.49 1062.0699 L921.31 1041.76 Z"
      /><path d="M921.31 1041.76 L948.85 1052.3199 L952 1080 L900.1 1080 L900.49 1062.0699 L921.31 1041.76 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M409.03 410.13 L427.16 428.26 L415.99 459.54 L383.32 456.18 L378.52 423 L409.03 410.13 Z"
      /><path d="M409.03 410.13 L427.16 428.26 L415.99 459.54 L383.32 456.18 L378.52 423 L409.03 410.13 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M951.84 632.89 L935.63 649.14 L949.66 684.81 L991.48 681.3 L993.99 670.18 L971.75 633.14 L951.84 632.89 Z"
      /><path d="M951.84 632.89 L935.63 649.14 L949.66 684.81 L991.48 681.3 L993.99 670.18 L971.75 633.14 L951.84 632.89 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1075.4301 927.39 L1061.53 926.05 L1035.45 961.97 L1042.24 976.05 L1072.5601 985.78 L1090.62 969.22 L1091.21 945.14 L1075.4301 927.39 Z"
      /><path d="M1075.4301 927.39 L1061.53 926.05 L1035.45 961.97 L1042.24 976.05 L1072.5601 985.78 L1090.62 969.22 L1091.21 945.14 L1075.4301 927.39 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1601.11 908.48 L1625.61 910.04 L1641.1899 955.33 L1619.58 968.91 L1580.3 948.58 L1576.95 937.25 L1601.11 908.48 Z"
      /><path d="M1601.11 908.48 L1625.61 910.04 L1641.1899 955.33 L1619.58 968.91 L1580.3 948.58 L1576.95 937.25 L1601.11 908.48 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M841.19 120.69 L817.12 89.61 L790.8 115.41 L795.5 129.14 L815.87 138.01 L841.19 120.69 Z"
      /><path d="M841.19 120.69 L817.12 89.61 L790.8 115.41 L795.5 129.14 L815.87 138.01 L841.19 120.69 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1641.37 235.61 L1654.2 246.08 L1650.98 275.8 L1610.75 284.8 L1601.08 257.8 L1615.63 237.32 L1641.37 235.61 Z"
      /><path d="M1641.37 235.61 L1654.2 246.08 L1650.98 275.8 L1610.75 284.8 L1601.08 257.8 L1615.63 237.32 L1641.37 235.61 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M431.39 167.69 L416.65 209.85 L453.62 230.51 L471.26 216.3 L470.27 187.93 L431.39 167.69 Z"
      /><path d="M431.39 167.69 L416.65 209.85 L453.62 230.51 L471.26 216.3 L470.27 187.93 L431.39 167.69 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1482.98 48.23 L1480.92 71.05 L1442.97 84.35 L1439.85 83.03 L1434.55 71.89 L1443.75 40.39 L1460.66 33.64 L1482.98 48.23 Z"
      /><path d="M1482.98 48.23 L1480.92 71.05 L1442.97 84.35 L1439.85 83.03 L1434.55 71.89 L1443.75 40.39 L1460.66 33.64 L1482.98 48.23 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M638.35 145.03 L621.14 154.44 L618.34 195.17 L642.48 212.11 L673.51 192.33 L674.77 157.64 L638.35 145.03 Z"
      /><path d="M638.35 145.03 L621.14 154.44 L618.34 195.17 L642.48 212.11 L673.51 192.33 L674.77 157.64 L638.35 145.03 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1167.66 33.83 L1180.3199 40.3 L1188.74 62.03 L1179.03 87.59 L1149.1801 78.26 L1139.11 53.82 L1142.02 45.85 L1167.66 33.83 Z"
      /><path d="M1167.66 33.83 L1180.3199 40.3 L1188.74 62.03 L1179.03 87.59 L1149.1801 78.26 L1139.11 53.82 L1142.02 45.85 L1167.66 33.83 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1901.87 49.45 L1885.8199 31.69 L1857.29 35.44 L1855.91 61.41 L1879.78 73.59 L1901.87 49.45 Z"
      /><path d="M1901.87 49.45 L1885.8199 31.69 L1857.29 35.44 L1855.91 61.41 L1879.78 73.59 L1901.87 49.45 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M383.32 456.18 L415.99 459.54 L426.41 474.82 L415.2 498.51 L379.93 504.84 L370.85 468.92 L383.32 456.18 Z"
      /><path d="M383.32 456.18 L415.99 459.54 L426.41 474.82 L415.2 498.51 L379.93 504.84 L370.85 468.92 L383.32 456.18 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M770.7 0 L815 0 L812.4 36.93 L781.96 35.92 L770.7 0 Z"
      /><path d="M770.7 0 L815 0 L812.4 36.93 L781.96 35.92 L770.7 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1258.97 556.57 L1274.72 568.38 L1277.6899 601.94 L1247.62 610.72 L1217.8199 582.09 L1229.52 563.84 L1258.97 556.57 Z"
      /><path d="M1258.97 556.57 L1274.72 568.38 L1277.6899 601.94 L1247.62 610.72 L1217.8199 582.09 L1229.52 563.84 L1258.97 556.57 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1773.99 253.27 L1755.76 250.33 L1736.47 270.39 L1747.03 305.42 L1774.54 302.74 L1786.64 275.57 L1773.99 253.27 Z"
      /><path d="M1773.99 253.27 L1755.76 250.33 L1736.47 270.39 L1747.03 305.42 L1774.54 302.74 L1786.64 275.57 L1773.99 253.27 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M873.76 551.83 L848.15 588.48 L879.82 612.59 L894.75 610.04 L906.46 596.44 L899.01 560.14 L873.76 551.83 Z"
      /><path d="M873.76 551.83 L848.15 588.48 L879.82 612.59 L894.75 610.04 L906.46 596.44 L899.01 560.14 L873.76 551.83 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M854.99 1045.95 L839.72 1034.54 L812.34 1044.52 L810.6 1080 L852.2 1080 L854.99 1045.95 Z"
      /><path d="M854.99 1045.95 L839.72 1034.54 L812.34 1044.52 L810.6 1080 L852.2 1080 L854.99 1045.95 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1080.6801 173.93 L1117.75 201.94 L1111.26 219.53 L1075.67 228.14 L1058.5 204.06 L1070.17 178.46 L1080.6801 173.93 Z"
      /><path d="M1080.6801 173.93 L1117.75 201.94 L1111.26 219.53 L1075.67 228.14 L1058.5 204.06 L1070.17 178.46 L1080.6801 173.93 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M359.82 987.3 L395.26 1009.09 L396.56 1027.0601 L376.77 1045.8199 L339.26 1030.47 L338.31 1008.3 L359.82 987.3 Z"
      /><path d="M359.82 987.3 L395.26 1009.09 L396.56 1027.0601 L376.77 1045.8199 L339.26 1030.47 L338.31 1008.3 L359.82 987.3 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1455.34 1052.53 L1420.17 1024.54 L1390.3199 1049.8101 L1389.8 1080 L1456.4 1080 L1455.34 1052.53 Z"
      /><path d="M1455.34 1052.53 L1420.17 1024.54 L1390.3199 1049.8101 L1389.8 1080 L1456.4 1080 L1455.34 1052.53 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1283.09 605.37 L1277.6899 601.94 L1247.62 610.72 L1236.6801 643.75 L1245.66 655.7 L1281.67 656.51 L1293.45 631.48 L1283.09 605.37 Z"
      /><path d="M1283.09 605.37 L1277.6899 601.94 L1247.62 610.72 L1236.6801 643.75 L1245.66 655.7 L1281.67 656.51 L1293.45 631.48 L1283.09 605.37 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1464.5 0 L1417.4 0 L1419.49 24.85 L1443.75 40.39 L1460.66 33.64 L1464.5 0 Z"
      /><path d="M1464.5 0 L1417.4 0 L1419.49 24.85 L1443.75 40.39 L1460.66 33.64 L1464.5 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1524.22 131.58 L1524.9301 148.16 L1498.1 173.88 L1492.88 174.36 L1478.36 159.64 L1492.3101 121.4 L1524.22 131.58 Z"
      /><path d="M1524.22 131.58 L1524.9301 148.16 L1498.1 173.88 L1492.88 174.36 L1478.36 159.64 L1492.3101 121.4 L1524.22 131.58 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M790.1 300.51 L752.9 269.91 L724.19 306.84 L764.33 336.19 L790.1 300.51 Z"
      /><path d="M790.1 300.51 L752.9 269.91 L724.19 306.84 L764.33 336.19 L790.1 300.51 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1814.84 921.49 L1837.64 936.51 L1842.27 962.59 L1825.72 978.93 L1792.24 976.03 L1775.95 952.44 L1777.9301 942.05 L1814.84 921.49 Z"
      /><path d="M1814.84 921.49 L1837.64 936.51 L1842.27 962.59 L1825.72 978.93 L1792.24 976.03 L1775.95 952.44 L1777.9301 942.05 L1814.84 921.49 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1871.04 788.85 L1857.22 787.4 L1830.84 815.43 L1836.8199 836.81 L1855.99 849.83 L1871.85 846.1 L1891.84 813.27 L1871.04 788.85 Z"
      /><path d="M1871.04 788.85 L1857.22 787.4 L1830.84 815.43 L1836.8199 836.81 L1855.99 849.83 L1871.85 846.1 L1891.84 813.27 L1871.04 788.85 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M253.93 89.53 L248.47 113.3 L209.93 112.07 L198.32 86.07 L231.27 63.19 L253.93 89.53 Z"
      /><path d="M253.93 89.53 L248.47 113.3 L209.93 112.07 L198.32 86.07 L231.27 63.19 L253.93 89.53 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M468.87 809.45 L454.1 795.44 L416.42 807.34 L411.99 829.27 L448.19 851.13 L465.8 839.93 L468.87 809.45 Z"
      /><path d="M468.87 809.45 L454.1 795.44 L416.42 807.34 L411.99 829.27 L448.19 851.13 L465.8 839.93 L468.87 809.45 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M999 744.52 L1014.68 747.47 L1032.83 779.36 L1019.72 803.99 L998.67 805.52 L976.48 776.41 L999 744.52 Z"
      /><path d="M999 744.52 L1014.68 747.47 L1032.83 779.36 L1019.72 803.99 L998.67 805.52 L976.48 776.41 L999 744.52 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M826.4 722.82 L787.64 733.54 L785.78 764.01 L820.74 773.07 L840.97 752.41 L826.4 722.82 Z"
      /><path d="M826.4 722.82 L787.64 733.54 L785.78 764.01 L820.74 773.07 L840.97 752.41 L826.4 722.82 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M656.77 554.38 L647.28 526.42 L608.37 528.57 L603.09 533.09 L605.78 571.7 L629.74 586.07 L639.38 583.65 L656.77 554.38 Z"
      /><path d="M656.77 554.38 L647.28 526.42 L608.37 528.57 L603.09 533.09 L605.78 571.7 L629.74 586.07 L639.38 583.65 L656.77 554.38 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M803.52 991.77 L793.69 1031.5 L772.72 1036.89 L753.92 1025.98 L752.37 1001.03 L775.3 981.35 L803.52 991.77 Z"
      /><path d="M803.52 991.77 L793.69 1031.5 L772.72 1036.89 L753.92 1025.98 L752.37 1001.03 L775.3 981.35 L803.52 991.77 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1392.8101 48.56 L1377.05 37.54 L1341.35 47.64 L1339.8101 69.47 L1349.85 82.34 L1382.79 83.73 L1395.3 58.58 L1392.8101 48.56 Z"
      /><path d="M1392.8101 48.56 L1377.05 37.54 L1341.35 47.64 L1339.8101 69.47 L1349.85 82.34 L1382.79 83.73 L1395.3 58.58 L1392.8101 48.56 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 137 L1920 178 L1883.54 184.29 L1858.49 144.87 L1858.49 144.85 L1863.37 138.52 L1920 137 Z"
      /><path d="M1920 137 L1920 178 L1883.54 184.29 L1858.49 144.87 L1858.49 144.85 L1863.37 138.52 L1920 137 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1692.26 288.19 L1710.03 315.54 L1693.98 342.71 L1680.03 345.36 L1656.22 320.97 L1665.37 291.54 L1692.26 288.19 Z"
      /><path d="M1692.26 288.19 L1710.03 315.54 L1693.98 342.71 L1680.03 345.36 L1656.22 320.97 L1665.37 291.54 L1692.26 288.19 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M407.4 0 L370 0 L368.56 52.99 L385.55 58.8 L415.19 47.05 L418.43 38.21 L407.4 0 Z"
      /><path d="M407.4 0 L370 0 L368.56 52.99 L385.55 58.8 L415.19 47.05 L418.43 38.21 L407.4 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1105.23 743.89 L1126.45 772.08 L1119.64 796.74 L1082.64 804.75 L1066.3 774.35 L1074 756.27 L1105.23 743.89 Z"
      /><path d="M1105.23 743.89 L1126.45 772.08 L1119.64 796.74 L1082.64 804.75 L1066.3 774.35 L1074 756.27 L1105.23 743.89 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1722.5699 367.48 L1719.8101 387.22 L1691.61 403.41 L1664.0699 374.41 L1680.03 345.36 L1693.98 342.71 L1722.5699 367.48 Z"
      /><path d="M1722.5699 367.48 L1719.8101 387.22 L1691.61 403.41 L1664.0699 374.41 L1680.03 345.36 L1693.98 342.71 L1722.5699 367.48 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M442.59 373.1 L442.7 373.13 L460.36 410.64 L453.87 424.48 L427.16 428.26 L409.03 410.13 L411.72 389.83 L442.59 373.1 Z"
      /><path d="M442.59 373.1 L442.7 373.13 L460.36 410.64 L453.87 424.48 L427.16 428.26 L409.03 410.13 L411.72 389.83 L442.59 373.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1189.52 834.64 L1173.15 810.06 L1135.65 816.87 L1129.64 844.87 L1143.17 861.32 L1183.55 849 L1189.52 834.64 Z"
      /><path d="M1189.52 834.64 L1173.15 810.06 L1135.65 816.87 L1129.64 844.87 L1143.17 861.32 L1183.55 849 L1189.52 834.64 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1464.64 445.41 L1435.39 412.23 L1407.6899 435.48 L1409.78 472.26 L1433.5699 482.78 L1462.55 464.68 L1464.64 445.41 Z"
      /><path d="M1464.64 445.41 L1435.39 412.23 L1407.6899 435.48 L1409.78 472.26 L1433.5699 482.78 L1462.55 464.68 L1464.64 445.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M789.71 401.09 L753.59 397.79 L737.98 427.65 L765.86 451.7 L786.23 442.63 L789.71 401.09 Z"
      /><path d="M789.71 401.09 L753.59 397.79 L737.98 427.65 L765.86 451.7 L786.23 442.63 L789.71 401.09 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M689.93 254.6 L644.06 234.27 L621.86 262.32 L654.94 298.62 L687.27 278.18 L689.93 254.6 Z"
      /><path d="M689.93 254.6 L644.06 234.27 L621.86 262.32 L654.94 298.62 L687.27 278.18 L689.93 254.6 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M720.91 307.45 L687.27 278.18 L654.94 298.62 L652.81 310.23 L677.15 338.2 L701.55 336.31 L720.91 307.45 Z"
      /><path d="M720.91 307.45 L687.27 278.18 L654.94 298.62 L652.81 310.23 L677.15 338.2 L701.55 336.31 L720.91 307.45 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1435.89 408.07 L1416.62 380.45 L1368.3 384.07 L1365.66 422.98 L1407.6899 435.48 L1435.39 412.23 L1435.89 408.07 Z"
      /><path d="M1435.89 408.07 L1416.62 380.45 L1368.3 384.07 L1365.66 422.98 L1407.6899 435.48 L1435.39 412.23 L1435.89 408.07 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M699.7 0 L743.3 0 L738.99 52.64 L733.4 55.09 L698.26 41.61 L699.7 0 Z"
      /><path d="M699.7 0 L743.3 0 L738.99 52.64 L733.4 55.09 L698.26 41.61 L699.7 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M425.28 339.7 L405.74 337.96 L385.1 362.8 L385.14 368.51 L411.72 389.83 L442.59 373.1 L425.28 339.7 Z"
      /><path d="M425.28 339.7 L405.74 337.96 L385.1 362.8 L385.14 368.51 L411.72 389.83 L442.59 373.1 L425.28 339.7 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M321.7 0 L266.9 0 L265.18 32.15 L292.32 56.26 L319.78 40.56 L321.7 0 Z"
      /><path d="M321.7 0 L266.9 0 L265.18 32.15 L292.32 56.26 L319.78 40.56 L321.7 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1860.83 255.88 L1873.87 264.45 L1876.25 296.22 L1839.52 307.88 L1829.85 301.92 L1821.96 276.34 L1829.28 262.87 L1860.83 255.88 Z"
      /><path d="M1860.83 255.88 L1873.87 264.45 L1876.25 296.22 L1839.52 307.88 L1829.85 301.92 L1821.96 276.34 L1829.28 262.87 L1860.83 255.88 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1662.66 573.54 L1694.01 590.7 L1694.23 600.99 L1669.3 622.55 L1647.49 615.53 L1644.1801 608.46 L1662.66 573.54 Z"
      /><path d="M1662.66 573.54 L1694.01 590.7 L1694.23 600.99 L1669.3 622.55 L1647.49 615.53 L1644.1801 608.46 L1662.66 573.54 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1496.15 670.39 L1469.23 661.89 L1448 687.18 L1483.0601 713.66 L1497.4399 704.62 L1496.15 670.39 Z"
      /><path d="M1496.15 670.39 L1469.23 661.89 L1448 687.18 L1483.0601 713.66 L1497.4399 704.62 L1496.15 670.39 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M72.11 871.41 L74.19 876.57 L29.07 914.03 L0 909.3 L0 850.8 L72.11 871.41 Z"
      /><path d="M72.11 871.41 L74.19 876.57 L29.07 914.03 L0 909.3 L0 850.8 L72.11 871.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M453.62 230.51 L451.17 250.84 L421.8 265.31 L397.99 245.7 L405.09 215.07 L416.65 209.85 L453.62 230.51 Z"
      /><path d="M453.62 230.51 L451.17 250.84 L421.8 265.31 L397.99 245.7 L405.09 215.07 L416.65 209.85 L453.62 230.51 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M0 267.8 L30.71 271.2 L36.19 290.19 L16.16 314.53 L0 315.1 L0 267.8 Z"
      /><path d="M0 267.8 L30.71 271.2 L36.19 290.19 L16.16 314.53 L0 315.1 L0 267.8 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1245.66 655.7 L1237.0699 690.06 L1259.28 711.73 L1287.9301 700.2 L1293.39 675.43 L1281.67 656.51 L1245.66 655.7 Z"
      /><path d="M1245.66 655.7 L1237.0699 690.06 L1259.28 711.73 L1287.9301 700.2 L1293.39 675.43 L1281.67 656.51 L1245.66 655.7 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1077.3199 612.16 L1110.45 612.58 L1125.02 634.37 L1102.67 667.12 L1069.74 649.45 L1077.3199 612.16 Z"
      /><path d="M1077.3199 612.16 L1110.45 612.58 L1125.02 634.37 L1102.67 667.12 L1069.74 649.45 L1077.3199 612.16 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1682.53 844.74 L1648.99 842.56 L1634.14 861.21 L1643.37 891.75 L1672.39 896.15 L1694.48 865.57 L1682.53 844.74 Z"
      /><path d="M1682.53 844.74 L1648.99 842.56 L1634.14 861.21 L1643.37 891.75 L1672.39 896.15 L1694.48 865.57 L1682.53 844.74 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1059.5 489.59 L1022.65 506.81 L1045.8 545.54 L1063.92 545.57 L1082.67 513.1 L1059.5 489.59 Z"
      /><path d="M1059.5 489.59 L1022.65 506.81 L1045.8 545.54 L1063.92 545.57 L1082.67 513.1 L1059.5 489.59 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M828.67 171.16 L820.51 165.31 L782.12 175.02 L781.08 195.16 L808.04 212.43 L832.42 199.33 L828.67 171.16 Z"
      /><path d="M828.67 171.16 L820.51 165.31 L782.12 175.02 L781.08 195.16 L808.04 212.43 L832.42 199.33 L828.67 171.16 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M465.8 839.93 L499.31 857.31 L485.5 893.6 L467.78 897.01 L443.67 875.98 L448.19 851.13 L465.8 839.93 Z"
      /><path d="M465.8 839.93 L499.31 857.31 L485.5 893.6 L467.78 897.01 L443.67 875.98 L448.19 851.13 L465.8 839.93 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M914.58 897.03 L897.3 889.54 L870.53 899.39 L863.13 916.03 L872.35 939.1 L914.2 944.68 L921.95 936.04 L914.58 897.03 Z"
      /><path d="M914.58 897.03 L897.3 889.54 L870.53 899.39 L863.13 916.03 L872.35 939.1 L914.2 944.68 L921.95 936.04 L914.58 897.03 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M587.31 746.73 L592.11 770.57 L561.24 794.95 L539.09 766.71 L550.55 738.73 L587.31 746.73 Z"
      /><path d="M587.31 746.73 L592.11 770.57 L561.24 794.95 L539.09 766.71 L550.55 738.73 L587.31 746.73 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1213.75 886.6 L1196.05 880.8 L1170.33 899.13 L1169.4 917.75 L1187.84 934.68 L1217.38 920.1 L1213.75 886.6 Z"
      /><path d="M1213.75 886.6 L1196.05 880.8 L1170.33 899.13 L1169.4 917.75 L1187.84 934.68 L1217.38 920.1 L1213.75 886.6 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1668.58 1021.83 L1684.42 1041.64 L1684.1 1080 L1601.6 1080 L1625.95 1023.34 L1668.58 1021.83 Z"
      /><path d="M1668.58 1021.83 L1684.42 1041.64 L1684.1 1080 L1601.6 1080 L1625.95 1023.34 L1668.58 1021.83 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1464.5 0 L1505.8 0 L1504.71 36.89 L1482.98 48.23 L1460.66 33.64 L1464.5 0 Z"
      /><path d="M1464.5 0 L1505.8 0 L1504.71 36.89 L1482.98 48.23 L1460.66 33.64 L1464.5 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1519.9399 468.17 L1492.12 488.01 L1491.87 506.53 L1509.62 522.51 L1544.47 515.82 L1547.08 479.64 L1519.9399 468.17 Z"
      /><path d="M1519.9399 468.17 L1492.12 488.01 L1491.87 506.53 L1509.62 522.51 L1544.47 515.82 L1547.08 479.64 L1519.9399 468.17 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M57.54 1043.71 L60.1 1080 L0 1080 L0 1050.3 L57.47 1043.63 L57.54 1043.71 Z"
      /><path d="M57.54 1043.71 L60.1 1080 L0 1080 L0 1050.3 L57.47 1043.63 L57.54 1043.71 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1063.92 545.57 L1045.8 545.54 L1024.35 567.74 L1040.74 599.75 L1068 601.08 L1080.29 565.58 L1063.92 545.57 Z"
      /><path d="M1063.92 545.57 L1045.8 545.54 L1024.35 567.74 L1040.74 599.75 L1068 601.08 L1080.29 565.58 L1063.92 545.57 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M1535.54 269.29 L1550.95 272.79 L1569.7 302.94 L1563.17 322.56 L1531.12 332.34 L1509.9 306.75 L1528.02 271.86 L1535.54 269.29 Z"
      /><path d="M1535.54 269.29 L1550.95 272.79 L1569.7 302.94 L1563.17 322.56 L1531.12 332.34 L1509.9 306.75 L1528.02 271.86 L1535.54 269.29 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M899.97 695.86 L937.27 703.97 L944.27 727.43 L937.77 740.62 L910.74 750.48 L885.39 735.96 L883.61 711.9 L899.97 695.86 Z"
      /><path d="M899.97 695.86 L937.27 703.97 L944.27 727.43 L937.77 740.62 L910.74 750.48 L885.39 735.96 L883.61 711.9 L899.97 695.86 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1827.46 631.28 L1863.5601 632.82 L1872.83 657.57 L1867.6 670.91 L1833.6801 681.29 L1812.64 651.51 L1827.46 631.28 Z"
      /><path d="M1827.46 631.28 L1863.5601 632.82 L1872.83 657.57 L1867.6 670.91 L1833.6801 681.29 L1812.64 651.51 L1827.46 631.28 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1375.6 0 L1417.4 0 L1419.49 24.85 L1392.8101 48.56 L1377.05 37.54 L1375.6 0 Z"
      /><path d="M1375.6 0 L1417.4 0 L1419.49 24.85 L1392.8101 48.56 L1377.05 37.54 L1375.6 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M945.38 879.16 L954.76 881.86 L971 913.61 L955.65 935.97 L921.95 936.04 L914.58 897.03 L945.38 879.16 Z"
      /><path d="M945.38 879.16 L954.76 881.86 L971 913.61 L955.65 935.97 L921.95 936.04 L914.58 897.03 L945.38 879.16 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M874.05 341.76 L895.63 356.02 L899.98 393.03 L877.75 406.2 L852.23 396.25 L847.78 361.89 L874.05 341.76 Z"
      /><path d="M874.05 341.76 L895.63 356.02 L899.98 393.03 L877.75 406.2 L852.23 396.25 L847.78 361.89 L874.05 341.76 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M177.13 47.26 L160.52 38.85 L134.03 52.18 L132.33 67.23 L159.05 96.42 L184.03 81.23 L177.13 47.26 Z"
      /><path d="M177.13 47.26 L160.52 38.85 L134.03 52.18 L132.33 67.23 L159.05 96.42 L184.03 81.23 L177.13 47.26 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1361.34 210.08 L1393.8199 217.74 L1403.2 235.67 L1378.1801 270.19 L1353.52 268.67 L1345.09 222.99 L1361.34 210.08 Z"
      /><path d="M1361.34 210.08 L1393.8199 217.74 L1403.2 235.67 L1378.1801 270.19 L1353.52 268.67 L1345.09 222.99 L1361.34 210.08 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M220.54 396.42 L236.9 414.18 L223.86 448.02 L183.79 442.98 L174.56 430.14 L195.57 396.47 L220.54 396.42 Z"
      /><path d="M220.54 396.42 L236.9 414.18 L223.86 448.02 L183.79 442.98 L174.56 430.14 L195.57 396.47 L220.54 396.42 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M285.58 371.81 L312.2 390.58 L311.67 414.39 L282.77 431.58 L259.37 411.88 L276.11 373.27 L285.58 371.81 Z"
      /><path d="M285.58 371.81 L312.2 390.58 L311.67 414.39 L282.77 431.58 L259.37 411.88 L276.11 373.27 L285.58 371.81 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M69.76 236.99 L56.14 252.55 L79.67 283.25 L92.69 281.25 L107.2 241.41 L106.32 239.18 L69.76 236.99 Z"
      /><path d="M69.76 236.99 L56.14 252.55 L79.67 283.25 L92.69 281.25 L107.2 241.41 L106.32 239.18 L69.76 236.99 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M233.15 359.58 L220.54 396.42 L195.57 396.47 L178.18 372.51 L185.14 350.2 L208.74 341.01 L233.15 359.58 Z"
      /><path d="M233.15 359.58 L220.54 396.42 L195.57 396.47 L178.18 372.51 L185.14 350.2 L208.74 341.01 L233.15 359.58 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M996.68 266.95 L977.87 248.46 L951.94 254.88 L941.73 271.16 L942.13 273.59 L970.15 296.5 L996.58 282.81 L996.68 266.95 Z"
      /><path d="M996.68 266.95 L977.87 248.46 L951.94 254.88 L941.73 271.16 L942.13 273.59 L970.15 296.5 L996.58 282.81 L996.68 266.95 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1574.97 573.44 L1550.25 559.79 L1530.1899 568.93 L1529.54 602.54 L1551.4 616.69 L1551.83 616.65 L1578.02 583.8 L1574.97 573.44 Z"
      /><path d="M1574.97 573.44 L1550.25 559.79 L1530.1899 568.93 L1529.54 602.54 L1551.4 616.69 L1551.83 616.65 L1578.02 583.8 L1574.97 573.44 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1396.53 160.83 L1412.03 185.89 L1393.8199 217.74 L1361.34 210.08 L1358.66 177.07 L1396.53 160.83 Z"
      /><path d="M1396.53 160.83 L1412.03 185.89 L1393.8199 217.74 L1361.34 210.08 L1358.66 177.07 L1396.53 160.83 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M73.08 32.67 L84.8 46.12 L81.71 62.36 L50.45 77.12 L45.49 75.91 L33.21 44.77 L39.5 36.03 L73.08 32.67 Z"
      /><path d="M73.08 32.67 L84.8 46.12 L81.71 62.36 L50.45 77.12 L45.49 75.91 L33.21 44.77 L39.5 36.03 L73.08 32.67 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1857.29 35.44 L1852.85 30.64 L1819.15 32.56 L1811.0699 45.68 L1834.02 74.78 L1855.91 61.41 L1857.29 35.44 Z"
      /><path d="M1857.29 35.44 L1852.85 30.64 L1819.15 32.56 L1811.0699 45.68 L1834.02 74.78 L1855.91 61.41 L1857.29 35.44 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 1080 L1861.1 1080 L1868.71 1046.59 L1920 1046.3 L1920 1080 Z"
      /><path d="M1920 1080 L1861.1 1080 L1868.71 1046.59 L1920 1046.3 L1920 1080 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1015.37 504.89 L1022.65 506.81 L1045.8 545.54 L1024.35 567.74 L1006.16 565.94 L989.06 530.77 L1015.37 504.89 Z"
      /><path d="M1015.37 504.89 L1022.65 506.81 L1045.8 545.54 L1024.35 567.74 L1006.16 565.94 L989.06 530.77 L1015.37 504.89 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M1739.49 850.18 L1780.6801 856.76 L1790.5699 868.77 L1790.62 869.19 L1756.72 909.05 L1735.35 904.98 L1721.8101 869.43 L1739.49 850.18 Z"
      /><path d="M1739.49 850.18 L1780.6801 856.76 L1790.5699 868.77 L1790.62 869.19 L1756.72 909.05 L1735.35 904.98 L1721.8101 869.43 L1739.49 850.18 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M117.22 954.11 L92.85 991.55 L61.1 992.87 L46.02 963.19 L51.16 949.59 L85.83 935.56 L117.22 954.11 Z"
      /><path d="M117.22 954.11 L92.85 991.55 L61.1 992.87 L46.02 963.19 L51.16 949.59 L85.83 935.56 L117.22 954.11 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1295.78 83.87 L1293.42 82.99 L1270.09 97.69 L1279 138.59 L1298.36 142.34 L1317.6899 119.5 L1295.78 83.87 Z"
      /><path d="M1295.78 83.87 L1293.42 82.99 L1270.09 97.69 L1279 138.59 L1298.36 142.34 L1317.6899 119.5 L1295.78 83.87 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1577.55 635.02 L1571.74 667.54 L1534.38 663.82 L1528.49 657.92 L1551.4 616.69 L1551.83 616.65 L1577.55 635.02 Z"
      /><path d="M1577.55 635.02 L1571.74 667.54 L1534.38 663.82 L1528.49 657.92 L1551.4 616.69 L1551.83 616.65 L1577.55 635.02 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M968.54 1031.25 L940.97 996.41 L917.04 1020.82 L921.31 1041.76 L948.85 1052.3199 L968.54 1031.25 Z"
      /><path d="M968.54 1031.25 L940.97 996.41 L917.04 1020.82 L921.31 1041.76 L948.85 1052.3199 L968.54 1031.25 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M873.73 333.95 L874.05 341.76 L847.78 361.89 L819.16 351.79 L820.14 307.27 L843.69 303.41 L873.73 333.95 Z"
      /><path d="M873.73 333.95 L874.05 341.76 L847.78 361.89 L819.16 351.79 L820.14 307.27 L843.69 303.41 L873.73 333.95 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1531.3101 51.27 L1504.71 36.89 L1482.98 48.23 L1480.92 71.05 L1495.9399 87.72 L1529.3199 80.05 L1531.3101 51.27 Z"
      /><path d="M1531.3101 51.27 L1504.71 36.89 L1482.98 48.23 L1480.92 71.05 L1495.9399 87.72 L1529.3199 80.05 L1531.3101 51.27 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M487.96 332.19 L520.45 351.88 L516.64 381.26 L501.86 390.47 L469.9 360.81 L479.87 334.79 L487.96 332.19 Z"
      /><path d="M487.96 332.19 L520.45 351.88 L516.64 381.26 L501.86 390.47 L469.9 360.81 L479.87 334.79 L487.96 332.19 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M103.2 624.55 L86.79 590.7 L50.04 595.43 L43.46 603.18 L56.62 654.41 L79.12 653.1 L103.2 624.55 Z"
      /><path d="M103.2 624.55 L86.79 590.7 L50.04 595.43 L43.46 603.18 L56.62 654.41 L79.12 653.1 L103.2 624.55 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M621.67 726.2 L644.56 755.74 L640.56 769.98 L617.67 783.67 L592.11 770.57 L587.31 746.73 L604.12 726.32 L621.67 726.2 Z"
      /><path d="M621.67 726.2 L644.56 755.74 L640.56 769.98 L617.67 783.67 L592.11 770.57 L587.31 746.73 L604.12 726.32 L621.67 726.2 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M158.14 99.31 L125.95 116.48 L122.77 131.98 L150.72 153.18 L171.68 131.44 L158.14 99.31 Z"
      /><path d="M158.14 99.31 L125.95 116.48 L122.77 131.98 L150.72 153.18 L171.68 131.44 L158.14 99.31 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1390.3199 1049.8101 L1357.4 1026.0601 L1333.4 1037.48 L1331.9 1080 L1389.8 1080 L1390.3199 1049.8101 Z"
      /><path d="M1390.3199 1049.8101 L1357.4 1026.0601 L1333.4 1037.48 L1331.9 1080 L1389.8 1080 L1390.3199 1049.8101 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1834.02 74.78 L1811.0699 45.68 L1787.1801 50.95 L1781.41 73.21 L1808.5 102.35 L1830.99 86.85 L1834.02 74.78 Z"
      /><path d="M1834.02 74.78 L1811.0699 45.68 L1787.1801 50.95 L1781.41 73.21 L1808.5 102.35 L1830.99 86.85 L1834.02 74.78 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1808.5 102.35 L1804.3199 118.91 L1797.21 125.32 L1740.98 103.56 L1746.4 89.11 L1781.41 73.21 L1808.5 102.35 Z"
      /><path d="M1808.5 102.35 L1804.3199 118.91 L1797.21 125.32 L1740.98 103.56 L1746.4 89.11 L1781.41 73.21 L1808.5 102.35 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1793.4399 323.28 L1774.54 302.74 L1747.03 305.42 L1740.16 313.65 L1748.77 351.56 L1766.85 357.8 L1793.33 339.37 L1793.4399 323.28 Z"
      /><path d="M1793.4399 323.28 L1774.54 302.74 L1747.03 305.42 L1740.16 313.65 L1748.77 351.56 L1766.85 357.8 L1793.33 339.37 L1793.4399 323.28 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M649.22 420.63 L619.77 429.11 L621.16 470.64 L639.61 476.76 L668.51 463.4 L666.46 433.01 L649.22 420.63 Z"
      /><path d="M649.22 420.63 L619.77 429.11 L621.16 470.64 L639.61 476.76 L668.51 463.4 L666.46 433.01 L649.22 420.63 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M712.24 461.71 L734.69 487.02 L732.37 495.31 L694.6 513.09 L686.54 509.02 L681.1 471.06 L712.24 461.71 Z"
      /><path d="M712.24 461.71 L734.69 487.02 L732.37 495.31 L694.6 513.09 L686.54 509.02 L681.1 471.06 L712.24 461.71 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1166.47 240.71 L1173.45 277.16 L1139.72 294.11 L1118.59 263.76 L1125.11 246.75 L1166.47 240.71 Z"
      /><path d="M1166.47 240.71 L1173.45 277.16 L1139.72 294.11 L1118.59 263.76 L1125.11 246.75 L1166.47 240.71 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M397.9 871.63 L418.35 886.73 L414.21 913.51 L372.15 919.63 L370.22 918.07 L367.83 885.59 L397.9 871.63 Z"
      /><path d="M397.9 871.63 L418.35 886.73 L414.21 913.51 L372.15 919.63 L370.22 918.07 L367.83 885.59 L397.9 871.63 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M512.72 915.98 L485.5 893.6 L467.78 897.01 L453.37 930.28 L469.39 952.48 L509.13 932.56 L512.72 915.98 Z"
      /><path d="M512.72 915.98 L485.5 893.6 L467.78 897.01 L453.37 930.28 L469.39 952.48 L509.13 932.56 L512.72 915.98 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1230.9 230.56 L1219.04 239.61 L1172.9 230.44 L1170.8 215.28 L1183.08 194.23 L1216.65 188.6 L1230.9 230.56 Z"
      /><path d="M1230.9 230.56 L1219.04 239.61 L1172.9 230.44 L1170.8 215.28 L1183.08 194.23 L1216.65 188.6 L1230.9 230.56 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M255.54 760.6 L209.29 730.02 L205.42 730.48 L187.8 771.72 L232.91 786.42 L253.71 770.18 L255.54 760.6 Z"
      /><path d="M255.54 760.6 L209.29 730.02 L205.42 730.48 L187.8 771.72 L232.91 786.42 L253.71 770.18 L255.54 760.6 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M891.19 231.55 L901.21 238.61 L904.99 256.18 L887.23 280.4 L861.05 276.9 L848.78 250.57 L854.45 240.71 L891.19 231.55 Z"
      /><path d="M891.19 231.55 L901.21 238.61 L904.99 256.18 L887.23 280.4 L861.05 276.9 L848.78 250.57 L854.45 240.71 L891.19 231.55 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1224.53 427.21 L1195.22 418.54 L1166.01 446.57 L1168.1899 467.78 L1193.79 478.96 L1222.38 464.89 L1224.53 427.21 Z"
      /><path d="M1224.53 427.21 L1195.22 418.54 L1166.01 446.57 L1168.1899 467.78 L1193.79 478.96 L1222.38 464.89 L1224.53 427.21 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M113.78 1034.2 L57.54 1043.71 L60.1 1080 L118.9 1080 L113.78 1034.2 Z"
      /><path d="M113.78 1034.2 L57.54 1043.71 L60.1 1080 L118.9 1080 L113.78 1034.2 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M407.4 0 L462.3 0 L458.44 25.86 L418.43 38.21 L407.4 0 Z"
      /><path d="M407.4 0 L462.3 0 L458.44 25.86 L418.43 38.21 L407.4 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M50.77 1012.27 L0 1008.5 L0 1050.3 L57.47 1043.63 L50.77 1012.27 Z"
      /><path d="M50.77 1012.27 L0 1008.5 L0 1050.3 L57.47 1043.63 L50.77 1012.27 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M314.73 906.87 L297.27 905.55 L270.79 931.66 L271.25 944.86 L302.93 965.68 L326.25 951.16 L330.59 926.39 L314.73 906.87 Z"
      /><path d="M314.73 906.87 L297.27 905.55 L270.79 931.66 L271.25 944.86 L302.93 965.68 L326.25 951.16 L330.59 926.39 L314.73 906.87 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M390.45 735.12 L359.56 738.1 L346.66 757.94 L364.81 789.89 L398.64 783.9 L407.52 758.11 L390.45 735.12 Z"
      /><path d="M390.45 735.12 L359.56 738.1 L346.66 757.94 L364.81 789.89 L398.64 783.9 L407.52 758.11 L390.45 735.12 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1395.3 58.58 L1382.79 83.73 L1392.8101 103.68 L1411.61 107.2 L1439.85 83.03 L1434.55 71.89 L1395.3 58.58 Z"
      /><path d="M1395.3 58.58 L1382.79 83.73 L1392.8101 103.68 L1411.61 107.2 L1439.85 83.03 L1434.55 71.89 L1395.3 58.58 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1428.64 619.02 L1398.9399 601.52 L1391.3 602.91 L1377.53 629.47 L1387.15 658.52 L1391.21 661.61 L1415.4399 656.69 L1431.4399 633.25 L1428.64 619.02 Z"
      /><path d="M1428.64 619.02 L1398.9399 601.52 L1391.3 602.91 L1377.53 629.47 L1387.15 658.52 L1391.21 661.61 L1415.4399 656.69 L1431.4399 633.25 L1428.64 619.02 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M735.51 111.62 L746.52 113.84 L760.31 156.27 L729.47 170.58 L706.89 148.93 L735.51 111.62 Z"
      /><path d="M735.51 111.62 L746.52 113.84 L760.31 156.27 L729.47 170.58 L706.89 148.93 L735.51 111.62 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1826.74 478.49 L1839.22 483.08 L1854.88 513.74 L1839.72 541.25 L1818.03 537.28 L1804.05 508.7 L1815.5601 483.61 L1826.74 478.49 Z"
      /><path d="M1826.74 478.49 L1839.22 483.08 L1854.88 513.74 L1839.72 541.25 L1818.03 537.28 L1804.05 508.7 L1815.5601 483.61 L1826.74 478.49 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M616.16 816.42 L610.85 821.19 L606.74 852.21 L627.41 869.85 L653.25 862.29 L660.31 827.04 L616.16 816.42 Z"
      /><path d="M616.16 816.42 L610.85 821.19 L606.74 852.21 L627.41 869.85 L653.25 862.29 L660.31 827.04 L616.16 816.42 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1527.38 747.7 L1490.74 756.74 L1488.4 763.71 L1502.21 798.77 L1510.1 802.19 L1535.9301 789.34 L1538.6899 757.67 L1527.38 747.7 Z"
      /><path d="M1527.38 747.7 L1490.74 756.74 L1488.4 763.71 L1502.21 798.77 L1510.1 802.19 L1535.9301 789.34 L1538.6899 757.67 L1527.38 747.7 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M686.63 745.43 L698.66 781.84 L671.18 799.59 L640.56 769.98 L644.56 755.74 L676.55 741.08 L686.63 745.43 Z"
      /><path d="M686.63 745.43 L698.66 781.84 L671.18 799.59 L640.56 769.98 L644.56 755.74 L676.55 741.08 L686.63 745.43 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1587.75 393.02 L1580.14 432.67 L1573.34 437.05 L1525.45 417.45 L1541.99 380.52 L1576.59 378.5 L1587.75 393.02 Z"
      /><path d="M1587.75 393.02 L1580.14 432.67 L1573.34 437.05 L1525.45 417.45 L1541.99 380.52 L1576.59 378.5 L1587.75 393.02 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1451.4 597.09 L1488.24 611.46 L1488.85 612.37 L1464.5601 645.32 L1431.4399 633.25 L1428.64 619.02 L1451.4 597.09 Z"
      /><path d="M1451.4 597.09 L1488.24 611.46 L1488.85 612.37 L1464.5601 645.32 L1431.4399 633.25 L1428.64 619.02 L1451.4 597.09 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1153.61 524.25 L1122.01 534.59 L1114.9399 563.27 L1126.53 579.04 L1151.22 582 L1173.71 558.86 L1172.95 535.64 L1153.61 524.25 Z"
      /><path d="M1153.61 524.25 L1122.01 534.59 L1114.9399 563.27 L1126.53 579.04 L1151.22 582 L1173.71 558.86 L1172.95 535.64 L1153.61 524.25 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1101.7 317.62 L1094.63 349.46 L1064.1 352.9 L1049.49 339.47 L1056.8 304.97 L1082.46 298.65 L1101.7 317.62 Z"
      /><path d="M1101.7 317.62 L1094.63 349.46 L1064.1 352.9 L1049.49 339.47 L1056.8 304.97 L1082.46 298.65 L1101.7 317.62 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1512.49 423.55 L1511.87 423.4 L1464.64 445.41 L1462.55 464.68 L1492.12 488.01 L1519.9399 468.17 L1512.49 423.55 Z"
      /><path d="M1512.49 423.55 L1511.87 423.4 L1464.64 445.41 L1462.55 464.68 L1492.12 488.01 L1519.9399 468.17 L1512.49 423.55 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M281.63 1007.9 L282.63 1030.8199 L256.47 1055.89 L219.85 1026.79 L219.29 1017.45 L246.3 991.33 L281.63 1007.9 Z"
      /><path d="M281.63 1007.9 L282.63 1030.8199 L256.47 1055.89 L219.85 1026.79 L219.29 1017.45 L246.3 991.33 L281.63 1007.9 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M858.82 652.73 L857.26 653.3 L847.69 697.79 L883.61 711.9 L899.97 695.86 L896.85 667.42 L858.82 652.73 Z"
      /><path d="M858.82 652.73 L857.26 653.3 L847.69 697.79 L883.61 711.9 L899.97 695.86 L896.85 667.42 L858.82 652.73 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M481.54 99.1 L466.61 62.62 L434.71 69.75 L428.61 101.91 L478.6 103.61 L481.54 99.1 Z"
      /><path d="M481.54 99.1 L466.61 62.62 L434.71 69.75 L428.61 101.91 L478.6 103.61 L481.54 99.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M748.15 526.47 L732.37 495.31 L694.6 513.09 L707.8 552.6 L717.06 553.07 L748.15 526.47 Z"
      /><path d="M748.15 526.47 L732.37 495.31 L694.6 513.09 L707.8 552.6 L717.06 553.07 L748.15 526.47 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M227.9 518.33 L250.79 526.44 L255.42 535.85 L246.97 573.41 L237.33 579.2 L197.79 565.9 L190.14 550.37 L191.45 545.43 L227.9 518.33 Z"
      /><path d="M227.9 518.33 L250.79 526.44 L255.42 535.85 L246.97 573.41 L237.33 579.2 L197.79 565.9 L190.14 550.37 L191.45 545.43 L227.9 518.33 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M116.8 0 L114.54 37.01 L134.03 52.18 L160.52 38.85 L157.7 0 L116.8 0 Z"
      /><path d="M116.8 0 L114.54 37.01 L134.03 52.18 L160.52 38.85 L157.7 0 L116.8 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M307.44 711.48 L308.05 751.12 L262.14 753.6 L264.03 719.36 L295.2 703.57 L307.44 711.48 Z"
      /><path d="M307.44 711.48 L308.05 751.12 L262.14 753.6 L264.03 719.36 L295.2 703.57 L307.44 711.48 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M434.71 69.75 L415.19 47.05 L385.55 58.8 L397.34 106.07 L424.42 105.93 L428.61 101.91 L434.71 69.75 Z"
      /><path d="M434.71 69.75 L415.19 47.05 L385.55 58.8 L397.34 106.07 L424.42 105.93 L428.61 101.91 L434.71 69.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1013.3 380.96 L1023.33 392.45 L1009.14 429.87 L979.53 429.52 L969.66 418.72 L975.92 380.31 L1013.3 380.96 Z"
      /><path d="M1013.3 380.96 L1023.33 392.45 L1009.14 429.87 L979.53 429.52 L969.66 418.72 L975.92 380.31 L1013.3 380.96 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1877.5601 452.64 L1874.15 467.04 L1839.22 483.08 L1826.74 478.49 L1828.1801 440.17 L1862.89 430.23 L1877.5601 452.64 Z"
      /><path d="M1877.5601 452.64 L1874.15 467.04 L1839.22 483.08 L1826.74 478.49 L1828.1801 440.17 L1862.89 430.23 L1877.5601 452.64 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M985.18 585.7 L991.33 612.93 L971.75 633.14 L951.84 632.89 L938.43 597.59 L955.04 577.23 L985.18 585.7 Z"
      /><path d="M985.18 585.7 L991.33 612.93 L971.75 633.14 L951.84 632.89 L938.43 597.59 L955.04 577.23 L985.18 585.7 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M706.89 148.93 L729.47 170.58 L726.75 198.67 L707.76 211.4 L673.51 192.33 L674.77 157.64 L689.01 147.67 L706.89 148.93 Z"
      /><path d="M706.89 148.93 L729.47 170.58 L726.75 198.67 L707.76 211.4 L673.51 192.33 L674.77 157.64 L689.01 147.67 L706.89 148.93 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1006.16 565.94 L1024.35 567.74 L1040.74 599.75 L1022.44 621.49 L991.33 612.93 L985.18 585.7 L1006.16 565.94 Z"
      /><path d="M1006.16 565.94 L1024.35 567.74 L1040.74 599.75 L1022.44 621.49 L991.33 612.93 L985.18 585.7 L1006.16 565.94 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M808.04 212.43 L781.08 195.16 L758.09 212.02 L762.93 247.53 L805.24 244.96 L808.04 212.43 Z"
      /><path d="M808.04 212.43 L781.08 195.16 L758.09 212.02 L762.93 247.53 L805.24 244.96 L808.04 212.43 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1149.99 483.05 L1117 478.95 L1099.58 511.37 L1122.01 534.59 L1153.61 524.25 L1149.99 483.05 Z"
      /><path d="M1149.99 483.05 L1117 478.95 L1099.58 511.37 L1122.01 534.59 L1153.61 524.25 L1149.99 483.05 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M163.42 709.4 L185.83 710.79 L205.42 730.48 L187.8 771.72 L183.51 774.17 L145.37 759.14 L143.18 728.36 L163.42 709.4 Z"
      /><path d="M163.42 709.4 L185.83 710.79 L205.42 730.48 L187.8 771.72 L183.51 774.17 L145.37 759.14 L143.18 728.36 L163.42 709.4 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M995.1 0 L954.6 0 L949.71 24.77 L975.05 56.27 L982.91 54.64 L1000.83 28.15 L995.1 0 Z"
      /><path d="M995.1 0 L954.6 0 L949.71 24.77 L975.05 56.27 L982.91 54.64 L1000.83 28.15 L995.1 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1230.9 230.56 L1242.95 231.69 L1264.74 269.07 L1246.76 290.96 L1213.51 275.7 L1219.04 239.61 L1230.9 230.56 Z"
      /><path d="M1230.9 230.56 L1242.95 231.69 L1264.74 269.07 L1246.76 290.96 L1213.51 275.7 L1219.04 239.61 L1230.9 230.56 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1529.54 602.54 L1495.33 614.46 L1516.9 656.49 L1528.49 657.92 L1551.4 616.69 L1529.54 602.54 Z"
      /><path d="M1529.54 602.54 L1495.33 614.46 L1516.9 656.49 L1528.49 657.92 L1551.4 616.69 L1529.54 602.54 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1705.99 265.71 L1692.26 288.19 L1710.03 315.54 L1740.16 313.65 L1747.03 305.42 L1736.47 270.39 L1705.99 265.71 Z"
      /><path d="M1705.99 265.71 L1692.26 288.19 L1710.03 315.54 L1740.16 313.65 L1747.03 305.42 L1736.47 270.39 L1705.99 265.71 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M0 447.1 L0 495.6 L48.21 496.29 L62.68 473.18 L52.48 449.94 L0 447.1 Z"
      /><path d="M0 447.1 L0 495.6 L48.21 496.29 L62.68 473.18 L52.48 449.94 L0 447.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1891.08 491.03 L1874.15 467.04 L1839.22 483.08 L1854.88 513.74 L1880.33 511.17 L1891.08 491.03 Z"
      /><path d="M1891.08 491.03 L1874.15 467.04 L1839.22 483.08 L1854.88 513.74 L1880.33 511.17 L1891.08 491.03 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M364.01 116.12 L342.59 90.3 L309.03 99.61 L305.2 114.94 L334.9 151.1 L335.66 150.99 L364.01 116.12 Z"
      /><path d="M364.01 116.12 L342.59 90.3 L309.03 99.61 L305.2 114.94 L334.9 151.1 L335.66 150.99 L364.01 116.12 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1143.17 861.32 L1129.64 844.87 L1092.49 851.62 L1084.63 868.16 L1100.0601 894.58 L1119.51 898.27 L1142.4 877.99 L1143.17 861.32 Z"
      /><path d="M1143.17 861.32 L1129.64 844.87 L1092.49 851.62 L1084.63 868.16 L1100.0601 894.58 L1119.51 898.27 L1142.4 877.99 L1143.17 861.32 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M251.75 355.45 L233.15 359.58 L220.54 396.42 L236.9 414.18 L259.37 411.88 L276.11 373.27 L251.75 355.45 Z"
      /><path d="M251.75 355.45 L233.15 359.58 L220.54 396.42 L236.9 414.18 L259.37 411.88 L276.11 373.27 L251.75 355.45 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1868.6801 595.2 L1839.35 584.36 L1817.36 597.22 L1827.46 631.28 L1863.5601 632.82 L1873.03 615.44 L1868.6801 595.2 Z"
      /><path d="M1868.6801 595.2 L1839.35 584.36 L1817.36 597.22 L1827.46 631.28 L1863.5601 632.82 L1873.03 615.44 L1868.6801 595.2 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1647.49 615.53 L1669.3 622.55 L1679.0699 648.03 L1668.29 660.2 L1640.3199 658.58 L1629.6899 647.33 L1647.49 615.53 Z"
      /><path d="M1647.49 615.53 L1669.3 622.55 L1679.0699 648.03 L1668.29 660.2 L1640.3199 658.58 L1629.6899 647.33 L1647.49 615.53 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1022.59 227.53 L985.66 219.24 L977.87 248.46 L996.68 266.95 L1027 245.77 L1022.59 227.53 Z"
      /><path d="M1022.59 227.53 L985.66 219.24 L977.87 248.46 L996.68 266.95 L1027 245.77 L1022.59 227.53 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M0 546.2 L37.91 550.47 L50.04 595.43 L43.46 603.18 L0 607.1 L0 546.2 Z"
      /><path d="M0 546.2 L37.91 550.47 L50.04 595.43 L43.46 603.18 L0 607.1 L0 546.2 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M63.02 421.69 L52.48 449.94 L0 447.1 L0 410.6 L43.42 401.24 L63.02 421.69 Z"
      /><path d="M63.02 421.69 L52.48 449.94 L0 447.1 L0 410.6 L43.42 401.24 L63.02 421.69 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1377.53 629.47 L1338.09 626.6 L1332.53 633.94 L1336.8101 668.87 L1337.3101 669.32 L1387.15 658.52 L1377.53 629.47 Z"
      /><path d="M1377.53 629.47 L1338.09 626.6 L1332.53 633.94 L1336.8101 668.87 L1337.3101 669.32 L1387.15 658.52 L1377.53 629.47 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 415.8 L1874.17 403.56 L1898.47 362.06 L1920 362 L1920 415.8 Z"
      /><path d="M1920 415.8 L1874.17 403.56 L1898.47 362.06 L1920 362 L1920 415.8 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1541.99 380.52 L1524.1899 355.32 L1482.1899 366.03 L1478.49 383.39 L1511.87 423.4 L1512.49 423.55 L1525.45 417.45 L1541.99 380.52 Z"
      /><path d="M1541.99 380.52 L1524.1899 355.32 L1482.1899 366.03 L1478.49 383.39 L1511.87 423.4 L1512.49 423.55 L1525.45 417.45 L1541.99 380.52 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1721.8101 869.43 L1694.48 865.57 L1672.39 896.15 L1686.6801 923.82 L1709.85 928.62 L1735.35 904.98 L1721.8101 869.43 Z"
      /><path d="M1721.8101 869.43 L1694.48 865.57 L1672.39 896.15 L1686.6801 923.82 L1709.85 928.62 L1735.35 904.98 L1721.8101 869.43 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1774.8101 388.99 L1809.42 397.88 L1810.09 425.14 L1774.8 446.52 L1750.6899 427.12 L1750.48 411.22 L1774.8101 388.99 Z"
      /><path d="M1774.8101 388.99 L1809.42 397.88 L1810.09 425.14 L1774.8 446.52 L1750.6899 427.12 L1750.48 411.22 L1774.8101 388.99 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1738.15 671.08 L1715.08 669.86 L1694.49 696.82 L1699.78 713.58 L1715.4399 722.56 L1739.62 713.88 L1746.17 679.46 L1738.15 671.08 Z"
      /><path d="M1738.15 671.08 L1715.08 669.86 L1694.49 696.82 L1699.78 713.58 L1715.4399 722.56 L1739.62 713.88 L1746.17 679.46 L1738.15 671.08 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1464.5601 645.32 L1431.4399 633.25 L1415.4399 656.69 L1443.29 688.24 L1448 687.18 L1469.23 661.89 L1464.5601 645.32 Z"
      /><path d="M1464.5601 645.32 L1431.4399 633.25 L1415.4399 656.69 L1443.29 688.24 L1448 687.18 L1469.23 661.89 L1464.5601 645.32 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1495.9399 87.72 L1480.92 71.05 L1442.97 84.35 L1458.88 114.22 L1488.72 115.82 L1495.9399 87.72 Z"
      /><path d="M1495.9399 87.72 L1480.92 71.05 L1442.97 84.35 L1458.88 114.22 L1488.72 115.82 L1495.9399 87.72 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M656.77 554.38 L696.49 561.95 L692.88 597.46 L669.86 606.61 L639.38 583.65 L656.77 554.38 Z"
      /><path d="M656.77 554.38 L696.49 561.95 L692.88 597.46 L669.86 606.61 L639.38 583.65 L656.77 554.38 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1126.39 1002.39 L1107.39 1018.21 L1107.83 1041.97 L1119.85 1053.75 L1153.55 1038.74 L1147.26 1010.64 L1126.39 1002.39 Z"
      /><path d="M1126.39 1002.39 L1107.39 1018.21 L1107.83 1041.97 L1119.85 1053.75 L1153.55 1038.74 L1147.26 1010.64 L1126.39 1002.39 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1307.8199 181.41 L1321.9 218.59 L1299.6 236.39 L1267.59 215.7 L1271.65 191.72 L1307.8199 181.41 Z"
      /><path d="M1307.8199 181.41 L1321.9 218.59 L1299.6 236.39 L1267.59 215.7 L1271.65 191.72 L1307.8199 181.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M988.16 727.94 L944.27 727.43 L937.77 740.62 L958.56 776.81 L976.48 776.41 L999 744.52 L988.16 727.94 Z"
      /><path d="M988.16 727.94 L944.27 727.43 L937.77 740.62 L958.56 776.81 L976.48 776.41 L999 744.52 L988.16 727.94 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M160.07 327.09 L132.36 340.13 L129.93 366.74 L142.69 381.18 L178.18 372.51 L185.14 350.2 L160.07 327.09 Z"
      /><path d="M160.07 327.09 L132.36 340.13 L129.93 366.74 L142.69 381.18 L178.18 372.51 L185.14 350.2 L160.07 327.09 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M694.6 513.09 L686.54 509.02 L650.16 522.05 L647.28 526.42 L656.77 554.38 L696.49 561.95 L707.8 552.6 L694.6 513.09 Z"
      /><path d="M694.6 513.09 L686.54 509.02 L650.16 522.05 L647.28 526.42 L656.77 554.38 L696.49 561.95 L707.8 552.6 L694.6 513.09 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M733.93 731.16 L740.71 762.95 L714.19 786.36 L698.66 781.84 L686.63 745.43 L724.43 726.1 L733.93 731.16 Z"
      /><path d="M733.93 731.16 L740.71 762.95 L714.19 786.36 L698.66 781.84 L686.63 745.43 L724.43 726.1 L733.93 731.16 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M594.02 945.59 L568.86 936.52 L551.47 959.1 L568.12 993.83 L606.17 977.75 L594.02 945.59 Z"
      /><path d="M594.02 945.59 L568.86 936.52 L551.47 959.1 L568.12 993.83 L606.17 977.75 L594.02 945.59 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1450.55 841.9 L1417.76 816.16 L1416.72 816.25 L1392.92 858.01 L1437.03 869.46 L1450.55 841.9 Z"
      /><path d="M1450.55 841.9 L1417.76 816.16 L1416.72 816.25 L1392.92 858.01 L1437.03 869.46 L1450.55 841.9 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1107.39 1018.21 L1107.83 1041.97 L1072.4 1052.15 L1057.84 1032.58 L1076.9301 1005.25 L1107.39 1018.21 Z"
      /><path d="M1107.39 1018.21 L1107.83 1041.97 L1072.4 1052.15 L1057.84 1032.58 L1076.9301 1005.25 L1107.39 1018.21 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M919.3 510.83 L919.85 546.25 L899.01 560.14 L873.76 551.83 L869.15 542.3 L887.61 501.45 L899.95 498.36 L919.3 510.83 Z"
      /><path d="M919.3 510.83 L919.85 546.25 L899.01 560.14 L873.76 551.83 L869.15 542.3 L887.61 501.45 L899.95 498.36 L919.3 510.83 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M1862.46 728.25 L1826.96 701.99 L1809.04 711.71 L1814.54 756.59 L1839.4 759.4 L1862.46 728.25 Z"
      /><path d="M1862.46 728.25 L1826.96 701.99 L1809.04 711.71 L1814.54 756.59 L1839.4 759.4 L1862.46 728.25 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M59.63 808.74 L0 825.7 L0 850.8 L72.11 871.41 L78.84 831.05 L59.63 808.74 Z"
      /><path d="M59.63 808.74 L0 825.7 L0 850.8 L72.11 871.41 L78.84 831.05 L59.63 808.74 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1630.79 391.64 L1637.89 423.52 L1616.85 443.42 L1580.14 432.67 L1587.75 393.02 L1630.79 391.64 Z"
      /><path d="M1630.79 391.64 L1637.89 423.52 L1616.85 443.42 L1580.14 432.67 L1587.75 393.02 L1630.79 391.64 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1584.99 770.94 L1614.12 771.64 L1620.66 807.62 L1600.45 820.23 L1568.92 806.78 L1584.99 770.94 Z"
      /><path d="M1584.99 770.94 L1614.12 771.64 L1620.66 807.62 L1600.45 820.23 L1568.92 806.78 L1584.99 770.94 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1524.9301 148.16 L1550.15 170.6 L1529.48 194.77 L1498.1 173.88 L1524.9301 148.16 Z"
      /><path d="M1524.9301 148.16 L1550.15 170.6 L1529.48 194.77 L1498.1 173.88 L1524.9301 148.16 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M959.34 161.09 L943.1 152.5 L916.46 167.32 L913.66 187.04 L939.74 209.75 L939.82 209.71 L962.25 174.19 L959.34 161.09 Z"
      /><path d="M959.34 161.09 L943.1 152.5 L916.46 167.32 L913.66 187.04 L939.74 209.75 L939.82 209.71 L962.25 174.19 L959.34 161.09 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1839.72 541.25 L1818.03 537.28 L1797.5601 554.74 L1799.21 591 L1817.36 597.22 L1839.35 584.36 L1841.55 543.97 L1839.72 541.25 Z"
      /><path d="M1839.72 541.25 L1818.03 537.28 L1797.5601 554.74 L1799.21 591 L1817.36 597.22 L1839.35 584.36 L1841.55 543.97 L1839.72 541.25 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M242.61 882.45 L237.46 906.55 L212.51 920.33 L183.95 902.17 L183.41 873.91 L213.95 853.95 L242.61 882.45 Z"
      /><path d="M242.61 882.45 L237.46 906.55 L212.51 920.33 L183.95 902.17 L183.41 873.91 L213.95 853.95 L242.61 882.45 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1049.77 448.68 L1024 447.36 L1005.05 483.78 L1015.37 504.89 L1022.65 506.81 L1059.5 489.59 L1063.16 463.82 L1049.77 448.68 Z"
      /><path d="M1049.77 448.68 L1024 447.36 L1005.05 483.78 L1015.37 504.89 L1022.65 506.81 L1059.5 489.59 L1063.16 463.82 L1049.77 448.68 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M848.15 588.48 L879.82 612.59 L858.82 652.73 L857.26 653.3 L833.53 643.96 L825.12 610.23 L842.95 589.17 L848.15 588.48 Z"
      /><path d="M848.15 588.48 L879.82 612.59 L858.82 652.73 L857.26 653.3 L833.53 643.96 L825.12 610.23 L842.95 589.17 L848.15 588.48 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1879.51 554.77 L1884.54 576.37 L1868.6801 595.2 L1839.35 584.36 L1841.55 543.97 L1879.51 554.77 Z"
      /><path d="M1879.51 554.77 L1884.54 576.37 L1868.6801 595.2 L1839.35 584.36 L1841.55 543.97 L1879.51 554.77 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 443.7 L1877.5601 452.64 L1874.15 467.04 L1891.08 491.03 L1920 488.6 L1920 443.7 Z"
      /><path d="M1920 443.7 L1877.5601 452.64 L1874.15 467.04 L1891.08 491.03 L1920 488.6 L1920 443.7 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M900.09 794.63 L872.13 789.82 L850.42 810.78 L864.87 842.26 L894.98 844.17 L900.52 839.99 L900.09 794.63 Z"
      /><path d="M900.09 794.63 L872.13 789.82 L850.42 810.78 L864.87 842.26 L894.98 844.17 L900.52 839.99 L900.09 794.63 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M565.97 999.27 L576.56 1028.41 L565.94 1043 L527.33 1043 L519.06 1032.0601 L524.32 1007.81 L565.97 999.27 Z"
      /><path d="M565.97 999.27 L576.56 1028.41 L565.94 1043 L527.33 1043 L519.06 1032.0601 L524.32 1007.81 L565.97 999.27 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M409.87 960.75 L379.2 954.88 L359.87 974.15 L359.82 987.3 L395.26 1009.09 L421.14 981.81 L409.87 960.75 Z"
      /><path d="M409.87 960.75 L379.2 954.88 L359.87 974.15 L359.82 987.3 L395.26 1009.09 L421.14 981.81 L409.87 960.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M615.46 263.35 L590.12 305.37 L582.98 305.27 L549.22 275.88 L549.14 273.54 L579.02 240.46 L615.46 263.35 Z"
      /><path d="M615.46 263.35 L590.12 305.37 L582.98 305.27 L549.22 275.88 L549.14 273.54 L579.02 240.46 L615.46 263.35 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M603.09 533.09 L576.22 530.26 L549.36 553.89 L575.72 585.44 L605.78 571.7 L603.09 533.09 Z"
      /><path d="M603.09 533.09 L576.22 530.26 L549.36 553.89 L575.72 585.44 L605.78 571.7 L603.09 533.09 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1386.1801 326.64 L1424.74 348.3 L1416.62 380.45 L1368.3 384.07 L1367.0601 382.52 L1370.6801 333.49 L1386.1801 326.64 Z"
      /><path d="M1386.1801 326.64 L1424.74 348.3 L1416.62 380.45 L1368.3 384.07 L1367.0601 382.52 L1370.6801 333.49 L1386.1801 326.64 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M432.78 984.26 L421.14 981.81 L395.26 1009.09 L396.56 1027.0601 L429.65 1042 L457.29 1019.99 L432.78 984.26 Z"
      /><path d="M432.78 984.26 L421.14 981.81 L395.26 1009.09 L396.56 1027.0601 L429.65 1042 L457.29 1019.99 L432.78 984.26 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M653.25 862.29 L627.41 869.85 L618.61 902.53 L627.75 918.29 L629.93 919.28 L671.4 904.58 L674.67 881.7 L653.25 862.29 Z"
      /><path d="M653.25 862.29 L627.41 869.85 L618.61 902.53 L627.75 918.29 L629.93 919.28 L671.4 904.58 L674.67 881.7 L653.25 862.29 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1311.9 720.43 L1310.14 750.49 L1277.4301 760.51 L1254.46 734.96 L1259.28 711.73 L1287.9301 700.2 L1311.9 720.43 Z"
      /><path d="M1311.9 720.43 L1310.14 750.49 L1277.4301 760.51 L1254.46 734.96 L1259.28 711.73 L1287.9301 700.2 L1311.9 720.43 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1528.49 657.92 L1516.9 656.49 L1496.15 670.39 L1497.4399 704.62 L1528.27 713.07 L1534.63 708.33 L1534.38 663.82 L1528.49 657.92 Z"
      /><path d="M1528.49 657.92 L1516.9 656.49 L1496.15 670.39 L1497.4399 704.62 L1528.27 713.07 L1534.63 708.33 L1534.38 663.82 L1528.49 657.92 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1391.21 661.61 L1387.15 658.52 L1337.3101 669.32 L1344.97 703.61 L1353.65 708.31 L1389.28 691.76 L1391.21 661.61 Z"
      /><path d="M1391.21 661.61 L1387.15 658.52 L1337.3101 669.32 L1344.97 703.61 L1353.65 708.31 L1389.28 691.76 L1391.21 661.61 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1264.6 1080 L1239.04 1036.76 L1211.77 1047.34 L1209 1080 L1264.6 1080 Z"
      /><path d="M1264.6 1080 L1239.04 1036.76 L1211.77 1047.34 L1209 1080 L1264.6 1080 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1114.9399 563.27 L1126.53 579.04 L1110.45 612.58 L1077.3199 612.16 L1068 601.08 L1080.29 565.58 L1114.9399 563.27 Z"
      /><path d="M1114.9399 563.27 L1126.53 579.04 L1110.45 612.58 L1077.3199 612.16 L1068 601.08 L1080.29 565.58 L1114.9399 563.27 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M859.86 756.17 L840.97 752.41 L820.74 773.07 L826.61 806.98 L850.42 810.78 L872.13 789.82 L859.86 756.17 Z"
      /><path d="M859.86 756.17 L840.97 752.41 L820.74 773.07 L826.61 806.98 L850.42 810.78 L872.13 789.82 L859.86 756.17 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M223.86 448.02 L232.17 464.38 L217.6 490.94 L173.17 487.85 L183.79 442.98 L223.86 448.02 Z"
      /><path d="M223.86 448.02 L232.17 464.38 L217.6 490.94 L173.17 487.85 L183.79 442.98 L223.86 448.02 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1691.61 403.41 L1664.0699 374.41 L1639.16 379.22 L1630.79 391.64 L1637.89 423.52 L1671.58 435.08 L1687 425.41 L1691.61 403.41 Z"
      /><path d="M1691.61 403.41 L1664.0699 374.41 L1639.16 379.22 L1630.79 391.64 L1637.89 423.52 L1671.58 435.08 L1687 425.41 L1691.61 403.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M492.8 754.37 L455.54 767.65 L454.1 795.44 L468.87 809.45 L503.09 801.13 L508.48 772.43 L492.8 754.37 Z"
      /><path d="M492.8 754.37 L455.54 767.65 L454.1 795.44 L468.87 809.45 L503.09 801.13 L508.48 772.43 L492.8 754.37 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1485.6801 850.72 L1466.95 836.74 L1450.55 841.9 L1437.03 869.46 L1446.63 892.37 L1486.61 875.81 L1485.6801 850.72 Z"
      /><path d="M1485.6801 850.72 L1466.95 836.74 L1450.55 841.9 L1437.03 869.46 L1446.63 892.37 L1486.61 875.81 L1485.6801 850.72 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1149.1801 78.26 L1139.11 53.82 L1106.1 63.62 L1106.1 96.92 L1125.02 103.95 L1149.1801 78.26 Z"
      /><path d="M1149.1801 78.26 L1139.11 53.82 L1106.1 63.62 L1106.1 96.92 L1125.02 103.95 L1149.1801 78.26 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1528.02 271.86 L1492.97 250.46 L1479.9301 255.26 L1466.98 279.68 L1488.3101 307.47 L1509.9 306.75 L1528.02 271.86 Z"
      /><path d="M1528.02 271.86 L1492.97 250.46 L1479.9301 255.26 L1466.98 279.68 L1488.3101 307.47 L1509.9 306.75 L1528.02 271.86 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M677.15 338.2 L652.81 310.23 L617.62 331.02 L636.76 371.08 L654.49 377.03 L658.12 375.55 L677.15 338.2 Z"
      /><path d="M677.15 338.2 L652.81 310.23 L617.62 331.02 L636.76 371.08 L654.49 377.03 L658.12 375.55 L677.15 338.2 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1883.78 92.87 L1865.0699 111.69 L1863.37 138.52 L1920 137 L1920 102 L1883.78 92.87 Z"
      /><path d="M1883.78 92.87 L1865.0699 111.69 L1863.37 138.52 L1920 137 L1920 102 L1883.78 92.87 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1142.02 45.85 L1119.75 16.6 L1087.9301 40.84 L1086.89 48.06 L1106.1 63.62 L1139.11 53.82 L1142.02 45.85 Z"
      /><path d="M1142.02 45.85 L1119.75 16.6 L1087.9301 40.84 L1086.89 48.06 L1106.1 63.62 L1139.11 53.82 L1142.02 45.85 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1565.23 469.67 L1598.05 491.93 L1587.55 521.9 L1553.4399 524.47 L1544.47 515.82 L1547.08 479.64 L1565.23 469.67 Z"
      /><path d="M1565.23 469.67 L1598.05 491.93 L1587.55 521.9 L1553.4399 524.47 L1544.47 515.82 L1547.08 479.64 L1565.23 469.67 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M471.26 216.3 L512.13 230.52 L512.95 244.17 L486.14 275.55 L474.37 275.04 L451.17 250.84 L453.62 230.51 L471.26 216.3 Z"
      /><path d="M471.26 216.3 L512.13 230.52 L512.95 244.17 L486.14 275.55 L474.37 275.04 L451.17 250.84 L453.62 230.51 L471.26 216.3 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M230.73 824.75 L216.95 835.55 L213.95 853.95 L242.61 882.45 L275.64 869.04 L280.97 856.45 L267.97 830.51 L230.73 824.75 Z"
      /><path d="M230.73 824.75 L216.95 835.55 L213.95 853.95 L242.61 882.45 L275.64 869.04 L280.97 856.45 L267.97 830.51 L230.73 824.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1584.61 79.64 L1630.3101 95.66 L1631.48 99.71 L1612.4301 132.81 L1579.45 126.72 L1578.48 86.3 L1584.61 79.64 Z"
      /><path d="M1584.61 79.64 L1630.3101 95.66 L1631.48 99.71 L1612.4301 132.81 L1579.45 126.72 L1578.48 86.3 L1584.61 79.64 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M157.7 0 L160.52 38.85 L177.13 47.26 L209.56 30.24 L210 0 L157.7 0 Z"
      /><path d="M157.7 0 L160.52 38.85 L177.13 47.26 L209.56 30.24 L210 0 L157.7 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1750.6899 427.12 L1774.8 446.52 L1776.02 461.75 L1757.36 485.75 L1719.91 482.23 L1720.6801 445.89 L1750.6899 427.12 Z"
      /><path d="M1750.6899 427.12 L1774.8 446.52 L1776.02 461.75 L1757.36 485.75 L1719.91 482.23 L1720.6801 445.89 L1750.6899 427.12 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M735.51 111.62 L706.89 148.93 L689.01 147.67 L681.12 97.42 L683.79 94.77 L721.06 94.31 L735.51 111.62 Z"
      /><path d="M735.51 111.62 L706.89 148.93 L689.01 147.67 L681.12 97.42 L683.79 94.77 L721.06 94.31 L735.51 111.62 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M861.92 111.23 L893.5 134.16 L891.65 146.96 L869.9 161.34 L857.65 157.14 L845.53 121.23 L861.92 111.23 Z"
      /><path d="M861.92 111.23 L893.5 134.16 L891.65 146.96 L869.9 161.34 L857.65 157.14 L845.53 121.23 L861.92 111.23 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1597.6 1080 L1552.96 1018.15 L1520.9301 1038.36 L1520.3 1080 L1597.6 1080 Z"
      /><path d="M1597.6 1080 L1552.96 1018.15 L1520.9301 1038.36 L1520.3 1080 L1597.6 1080 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1279 138.59 L1298.36 142.34 L1312.6 172.23 L1307.8199 181.41 L1271.65 191.72 L1253.75 172.39 L1258.83 150.29 L1279 138.59 Z"
      /><path d="M1279 138.59 L1298.36 142.34 L1312.6 172.23 L1307.8199 181.41 L1271.65 191.72 L1253.75 172.39 L1258.83 150.29 L1279 138.59 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1338.7 0 L1293.8 0 L1298.71 36.45 L1334.9301 39.94 L1338.7 0 Z"
      /><path d="M1338.7 0 L1293.8 0 L1298.71 36.45 L1334.9301 39.94 L1338.7 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M364.01 116.12 L335.66 150.99 L372.08 175.33 L394.2 157.52 L383.97 117.24 L364.01 116.12 Z"
      /><path d="M364.01 116.12 L335.66 150.99 L372.08 175.33 L394.2 157.52 L383.97 117.24 L364.01 116.12 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1815.33 354.62 L1793.33 339.37 L1766.85 357.8 L1774.8101 388.99 L1809.42 397.88 L1811.33 396.03 L1815.33 354.62 Z"
      /><path d="M1815.33 354.62 L1793.33 339.37 L1766.85 357.8 L1774.8101 388.99 L1809.42 397.88 L1811.33 396.03 L1815.33 354.62 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M857.65 157.14 L828.67 171.16 L832.42 199.33 L845.03 205.61 L875.55 191.79 L869.9 161.34 L857.65 157.14 Z"
      /><path d="M857.65 157.14 L828.67 171.16 L832.42 199.33 L845.03 205.61 L875.55 191.79 L869.9 161.34 L857.65 157.14 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1612.4301 132.81 L1620.46 151.82 L1611.35 170.9 L1569.9 171.75 L1566.74 168.99 L1572.36 132.14 L1579.45 126.72 L1612.4301 132.81 Z"
      /><path d="M1612.4301 132.81 L1620.46 151.82 L1611.35 170.9 L1569.9 171.75 L1566.74 168.99 L1572.36 132.14 L1579.45 126.72 L1612.4301 132.81 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1036.8101 1031.1899 L1016.5 1080 L1069.2 1080 L1072.4 1052.15 L1057.84 1032.58 L1036.8101 1031.1899 Z"
      /><path d="M1036.8101 1031.1899 L1016.5 1080 L1069.2 1080 L1072.4 1052.15 L1057.84 1032.58 L1036.8101 1031.1899 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M707.8 552.6 L717.06 553.07 L746.56 582.18 L735.31 609.58 L718.37 614.82 L692.88 597.46 L696.49 561.95 L707.8 552.6 Z"
      /><path d="M707.8 552.6 L717.06 553.07 L746.56 582.18 L735.31 609.58 L718.37 614.82 L692.88 597.46 L696.49 561.95 L707.8 552.6 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M512.95 244.17 L549.14 273.54 L549.22 275.88 L526.15 301.36 L504.94 301.01 L486.14 275.55 L512.95 244.17 Z"
      /><path d="M512.95 244.17 L549.14 273.54 L549.22 275.88 L526.15 301.36 L504.94 301.01 L486.14 275.55 L512.95 244.17 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M875.24 1040.15 L900.49 1062.0699 L900.1 1080 L852.2 1080 L854.99 1045.95 L875.24 1040.15 Z"
      /><path d="M875.24 1040.15 L900.49 1062.0699 L900.1 1080 L852.2 1080 L854.99 1045.95 L875.24 1040.15 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1106.1 63.62 L1086.89 48.06 L1063.12 62.24 L1063.17 84.42 L1091.0601 103.39 L1106.1 96.92 L1106.1 63.62 Z"
      /><path d="M1106.1 63.62 L1086.89 48.06 L1063.12 62.24 L1063.17 84.42 L1091.0601 103.39 L1106.1 96.92 L1106.1 63.62 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1297.21 266.75 L1264.74 269.07 L1246.76 290.96 L1250.73 314.49 L1269.7 324.31 L1300.3101 306.44 L1300.01 269.75 L1297.21 266.75 Z"
      /><path d="M1297.21 266.75 L1264.74 269.07 L1246.76 290.96 L1250.73 314.49 L1269.7 324.31 L1300.3101 306.44 L1300.01 269.75 L1297.21 266.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1760.2 541.89 L1797.5601 554.74 L1799.21 591 L1787.78 596.18 L1748.92 579.08 L1760.2 541.89 Z"
      /><path d="M1760.2 541.89 L1797.5601 554.74 L1799.21 591 L1787.78 596.18 L1748.92 579.08 L1760.2 541.89 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1759.08 800.59 L1732.9301 817.04 L1739.49 850.18 L1780.6801 856.76 L1785.6899 810.85 L1759.08 800.59 Z"
      /><path d="M1759.08 800.59 L1732.9301 817.04 L1739.49 850.18 L1780.6801 856.76 L1785.6899 810.85 L1759.08 800.59 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 242.1 L1871.84 207.17 L1859.64 212.79 L1860.83 255.88 L1873.87 264.45 L1920 242.7 L1920 242.1 Z"
      /><path d="M1920 242.1 L1871.84 207.17 L1859.64 212.79 L1860.83 255.88 L1873.87 264.45 L1920 242.7 L1920 242.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M65.86 319.78 L38.53 333.85 L35.38 359.87 L47.09 371.1 L80.6 363.28 L83.7 334.45 L65.86 319.78 Z"
      /><path d="M65.86 319.78 L38.53 333.85 L35.38 359.87 L47.09 371.1 L80.6 363.28 L83.7 334.45 L65.86 319.78 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1799.21 591 L1787.78 596.18 L1773.97 629.96 L1793.23 652.88 L1812.64 651.51 L1827.46 631.28 L1817.36 597.22 L1799.21 591 Z"
      /><path d="M1799.21 591 L1787.78 596.18 L1773.97 629.96 L1793.23 652.88 L1812.64 651.51 L1827.46 631.28 L1817.36 597.22 L1799.21 591 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M851.97 34.74 L861.76 43.84 L850.02 73.53 L817.93 78.12 L815.99 75.57 L815.66 40.29 L851.97 34.74 Z"
      /><path d="M851.97 34.74 L861.76 43.84 L850.02 73.53 L817.93 78.12 L815.99 75.57 L815.66 40.29 L851.97 34.74 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M989.56 116.82 L971.65 107.1 L950.05 111.25 L937.75 128.48 L943.1 152.5 L959.34 161.09 L985.09 143.44 L990.54 119.73 L989.56 116.82 Z"
      /><path d="M989.56 116.82 L971.65 107.1 L950.05 111.25 L937.75 128.48 L943.1 152.5 L959.34 161.09 L985.09 143.44 L990.54 119.73 L989.56 116.82 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M738.98 372.29 L753.59 397.79 L737.98 427.65 L719.69 431.88 L700.52 417.35 L698.43 391.7 L721.04 370.37 L738.98 372.29 Z"
      /><path d="M738.98 372.29 L753.59 397.79 L737.98 427.65 L719.69 431.88 L700.52 417.35 L698.43 391.7 L721.04 370.37 L738.98 372.29 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M325.12 653.07 L347.75 691.29 L342.34 701.86 L307.44 711.48 L295.2 703.57 L289.8 681.11 L305.94 656.28 L325.12 653.07 Z"
      /><path d="M325.12 653.07 L347.75 691.29 L342.34 701.86 L307.44 711.48 L295.2 703.57 L289.8 681.11 L305.94 656.28 L325.12 653.07 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M92.69 281.25 L114.08 297.04 L111.6 323.27 L83.7 334.45 L65.86 319.78 L64.57 301.08 L79.67 283.25 L92.69 281.25 Z"
      /><path d="M92.69 281.25 L114.08 297.04 L111.6 323.27 L83.7 334.45 L65.86 319.78 L64.57 301.08 L79.67 283.25 L92.69 281.25 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1629.6899 647.33 L1618.72 647.15 L1596.96 677.49 L1611.78 695.81 L1634.17 693.12 L1640.3199 658.58 L1629.6899 647.33 Z"
      /><path d="M1629.6899 647.33 L1618.72 647.15 L1596.96 677.49 L1611.78 695.81 L1634.17 693.12 L1640.3199 658.58 L1629.6899 647.33 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M583.07 897.17 L618.61 902.53 L627.75 918.29 L594.02 945.59 L568.86 936.52 L566.49 927.27 L583.07 897.17 Z"
      /><path d="M583.07 897.17 L618.61 902.53 L627.75 918.29 L594.02 945.59 L568.86 936.52 L566.49 927.27 L583.07 897.17 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M150.41 1017.44 L115.71 1030.67 L113.78 1034.2 L118.9 1080 L181.8 1080 L183.08 1066.5601 L150.41 1017.44 Z"
      /><path d="M150.41 1017.44 L115.71 1030.67 L113.78 1034.2 L118.9 1080 L181.8 1080 L183.08 1066.5601 L150.41 1017.44 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M825.12 610.23 L792.98 607.6 L775.54 633.3 L804.87 660.08 L833.53 643.96 L825.12 610.23 Z"
      /><path d="M825.12 610.23 L792.98 607.6 L775.54 633.3 L804.87 660.08 L833.53 643.96 L825.12 610.23 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1404.45 537.68 L1403.91 540.07 L1369.59 557.15 L1352.8101 547.97 L1344.66 515.81 L1380.76 501.69 L1404.45 537.68 Z"
      /><path d="M1404.45 537.68 L1403.91 540.07 L1369.59 557.15 L1352.8101 547.97 L1344.66 515.81 L1380.76 501.69 L1404.45 537.68 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1350.8 270.86 L1300.01 269.75 L1300.3101 306.44 L1330.4301 324.89 L1342.34 320.92 L1350.8 270.86 Z"
      /><path d="M1350.8 270.86 L1300.01 269.75 L1300.3101 306.44 L1330.4301 324.89 L1342.34 320.92 L1350.8 270.86 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M239.36 680.64 L209.42 666.77 L205.02 668.1 L185.83 710.79 L205.42 730.48 L209.29 730.02 L240.68 702.81 L239.36 680.64 Z"
      /><path d="M239.36 680.64 L209.42 666.77 L205.02 668.1 L185.83 710.79 L205.42 730.48 L209.29 730.02 L240.68 702.81 L239.36 680.64 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M645.09 952.92 L669.39 959.85 L676.72 978.29 L657.94 1003.58 L623.12 996.34 L615.33 981.56 L645.09 952.92 Z"
      /><path d="M645.09 952.92 L669.39 959.85 L676.72 978.29 L657.94 1003.58 L623.12 996.34 L615.33 981.56 L645.09 952.92 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1327 792.95 L1363.77 805.77 L1361.03 836.66 L1331.6 849.42 L1305.04 814.21 L1327 792.95 Z"
      /><path d="M1327 792.95 L1363.77 805.77 L1361.03 836.66 L1331.6 849.42 L1305.04 814.21 L1327 792.95 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M486.14 275.55 L474.37 275.04 L447.68 310.39 L448.01 312.51 L479.87 334.79 L487.96 332.19 L504.94 301.01 L486.14 275.55 Z"
      /><path d="M486.14 275.55 L474.37 275.04 L447.68 310.39 L448.01 312.51 L479.87 334.79 L487.96 332.19 L504.94 301.01 L486.14 275.55 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M292.32 56.26 L289.56 74.7 L253.93 89.53 L231.27 63.19 L231.98 51.27 L265.18 32.15 L292.32 56.26 Z"
      /><path d="M292.32 56.26 L289.56 74.7 L253.93 89.53 L231.27 63.19 L231.98 51.27 L265.18 32.15 L292.32 56.26 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M971 913.61 L955.65 935.97 L973.36 970.28 L981.79 972.02 L1011.13 953.43 L1003.63 913.93 L971 913.61 Z"
      /><path d="M971 913.61 L955.65 935.97 L973.36 970.28 L981.79 972.02 L1011.13 953.43 L1003.63 913.93 L971 913.61 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M345.55 869.3 L337.43 869.88 L314.73 906.87 L330.59 926.39 L370.22 918.07 L367.83 885.59 L345.55 869.3 Z"
      /><path d="M345.55 869.3 L337.43 869.88 L314.73 906.87 L330.59 926.39 L370.22 918.07 L367.83 885.59 L345.55 869.3 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1731.4 0 L1779.5 0 L1774.55 37.37 L1737.02 40.24 L1731.4 0 Z"
      /><path d="M1731.4 0 L1779.5 0 L1774.55 37.37 L1737.02 40.24 L1731.4 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1336.17 598.08 L1325.14 588.32 L1283.09 605.37 L1293.45 631.48 L1332.53 633.94 L1338.09 626.6 L1336.17 598.08 Z"
      /><path d="M1336.17 598.08 L1325.14 588.32 L1283.09 605.37 L1293.45 631.48 L1332.53 633.94 L1338.09 626.6 L1336.17 598.08 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M60.04 531.31 L81.57 536.16 L95.5 576.8 L86.79 590.7 L50.04 595.43 L37.91 550.47 L60.04 531.31 Z"
      /><path d="M60.04 531.31 L81.57 536.16 L95.5 576.8 L86.79 590.7 L50.04 595.43 L37.91 550.47 L60.04 531.31 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1458.88 114.22 L1488.72 115.82 L1492.3101 121.4 L1478.36 159.64 L1454.28 158.16 L1441.92 139.24 L1458.88 114.22 Z"
      /><path d="M1458.88 114.22 L1488.72 115.82 L1492.3101 121.4 L1478.36 159.64 L1454.28 158.16 L1441.92 139.24 L1458.88 114.22 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M989.06 530.77 L971.5 529.71 L949.33 557.48 L955.04 577.23 L985.18 585.7 L1006.16 565.94 L989.06 530.77 Z"
      /><path d="M989.06 530.77 L971.5 529.71 L949.33 557.48 L955.04 577.23 L985.18 585.7 L1006.16 565.94 L989.06 530.77 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M1765.0601 197.15 L1754.21 172.13 L1710.73 178.37 L1707.4 184.11 L1725.12 219.18 L1742.04 222.3 L1765.0601 197.15 Z"
      /><path d="M1765.0601 197.15 L1754.21 172.13 L1710.73 178.37 L1707.4 184.11 L1725.12 219.18 L1742.04 222.3 L1765.0601 197.15 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1194.4301 316.57 L1223.54 331.81 L1222.4399 364.42 L1187.45 375.94 L1167.84 336.93 L1194.4301 316.57 Z"
      /><path d="M1194.4301 316.57 L1223.54 331.81 L1222.4399 364.42 L1187.45 375.94 L1167.84 336.93 L1194.4301 316.57 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1305.04 814.21 L1331.6 849.42 L1324.15 871.89 L1308.4399 878.52 L1280.14 867.75 L1274.58 833.23 L1289.9 814.35 L1305.04 814.21 Z"
      /><path d="M1305.04 814.21 L1331.6 849.42 L1324.15 871.89 L1308.4399 878.52 L1280.14 867.75 L1274.58 833.23 L1289.9 814.35 L1305.04 814.21 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M629.74 586.07 L616.99 622.23 L593.45 627.44 L571.96 599.49 L575.72 585.44 L605.78 571.7 L629.74 586.07 Z"
      /><path d="M629.74 586.07 L616.99 622.23 L593.45 627.44 L571.96 599.49 L575.72 585.44 L605.78 571.7 L629.74 586.07 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M61.1 992.87 L46.02 963.19 L0 971.9 L0 1008.5 L50.77 1012.27 L61.1 992.87 Z"
      /><path d="M61.1 992.87 L46.02 963.19 L0 971.9 L0 1008.5 L50.77 1012.27 L61.1 992.87 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M33.21 44.77 L45.49 75.91 L24.94 91.28 L0 88 L0 46.1 L33.21 44.77 Z"
      /><path d="M33.21 44.77 L45.49 75.91 L24.94 91.28 L0 88 L0 46.1 L33.21 44.77 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M840.3 1008.58 L811.46 988.76 L803.52 991.77 L793.69 1031.5 L812.34 1044.52 L839.72 1034.54 L840.3 1008.58 Z"
      /><path d="M840.3 1008.58 L811.46 988.76 L803.52 991.77 L793.69 1031.5 L812.34 1044.52 L839.72 1034.54 L840.3 1008.58 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M321.7 0 L370 0 L368.56 52.99 L352.34 59.64 L319.78 40.56 L321.7 0 Z"
      /><path d="M321.7 0 L370 0 L368.56 52.99 L352.34 59.64 L319.78 40.56 L321.7 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1122.01 534.59 L1114.9399 563.27 L1080.29 565.58 L1063.92 545.57 L1082.67 513.1 L1099.58 511.37 L1122.01 534.59 Z"
      /><path d="M1122.01 534.59 L1114.9399 563.27 L1080.29 565.58 L1063.92 545.57 L1082.67 513.1 L1099.58 511.37 L1122.01 534.59 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M178.18 372.51 L142.69 381.18 L139.94 402.42 L160.69 427.88 L174.56 430.14 L195.57 396.47 L178.18 372.51 Z"
      /><path d="M178.18 372.51 L142.69 381.18 L139.94 402.42 L160.69 427.88 L174.56 430.14 L195.57 396.47 L178.18 372.51 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M162.79 246.69 L175.47 250.2 L191.06 273.87 L185.91 293.31 L164.2 303.86 L139.51 285.26 L142.03 261.28 L162.79 246.69 Z"
      /><path d="M162.79 246.69 L175.47 250.2 L191.06 273.87 L185.91 293.31 L164.2 303.86 L139.51 285.26 L142.03 261.28 L162.79 246.69 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M466.73 500.79 L441.53 533.45 L446.53 541.53 L486.4 551.71 L501.97 523.26 L487.61 501.21 L466.73 500.79 Z"
      /><path d="M466.73 500.79 L441.53 533.45 L446.53 541.53 L486.4 551.71 L501.97 523.26 L487.61 501.21 L466.73 500.79 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M121.39 882.91 L81 881.65 L85.83 935.56 L117.22 954.11 L118.72 953.85 L144.08 932.08 L145.41 926.94 L121.39 882.91 Z"
      /><path d="M121.39 882.91 L81 881.65 L85.83 935.56 L117.22 954.11 L118.72 953.85 L144.08 932.08 L145.41 926.94 L121.39 882.91 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1068.66 249.97 L1089.85 272.08 L1082.46 298.65 L1056.8 304.97 L1040.0699 291.49 L1045.0601 257.25 L1068.66 249.97 Z"
      /><path d="M1068.66 249.97 L1089.85 272.08 L1082.46 298.65 L1056.8 304.97 L1040.0699 291.49 L1045.0601 257.25 L1068.66 249.97 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1765.52 753.44 L1804.4301 763.91 L1801.16 803.13 L1785.6899 810.85 L1759.08 800.59 L1754.55 764.79 L1765.52 753.44 Z"
      /><path d="M1765.52 753.44 L1804.4301 763.91 L1801.16 803.13 L1785.6899 810.85 L1759.08 800.59 L1754.55 764.79 L1765.52 753.44 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1256.1 0 L1214.8 0 L1211.52 21.38 L1235.37 55.6 L1255.8 43.42 L1256.1 0 Z"
      /><path d="M1256.1 0 L1214.8 0 L1211.52 21.38 L1235.37 55.6 L1255.8 43.42 L1256.1 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M708.1 839.98 L713.54 865.6 L674.67 881.7 L653.25 862.29 L660.31 827.04 L666.53 822.38 L708.1 839.98 Z"
      /><path d="M708.1 839.98 L713.54 865.6 L674.67 881.7 L653.25 862.29 L660.31 827.04 L666.53 822.38 L708.1 839.98 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M481.39 689.46 L463.86 663.1 L434.33 670.95 L427.02 701.99 L446.42 718.75 L470.92 712.95 L481.39 689.46 Z"
      /><path d="M481.39 689.46 L463.86 663.1 L434.33 670.95 L427.02 701.99 L446.42 718.75 L470.92 712.95 L481.39 689.46 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1750.48 411.22 L1719.8101 387.22 L1691.61 403.41 L1687 425.41 L1720.6801 445.89 L1750.6899 427.12 L1750.48 411.22 Z"
      /><path d="M1750.48 411.22 L1719.8101 387.22 L1691.61 403.41 L1687 425.41 L1720.6801 445.89 L1750.6899 427.12 L1750.48 411.22 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M799.89 362.43 L765.19 342.03 L738.98 372.29 L753.59 397.79 L789.71 401.09 L795.81 396.68 L799.89 362.43 Z"
      /><path d="M799.89 362.43 L765.19 342.03 L738.98 372.29 L753.59 397.79 L789.71 401.09 L795.81 396.68 L799.89 362.43 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1720.6801 445.89 L1719.91 482.23 L1716.37 485.51 L1685.23 487.01 L1667.64 468.75 L1671.58 435.08 L1687 425.41 L1720.6801 445.89 Z"
      /><path d="M1720.6801 445.89 L1719.91 482.23 L1716.37 485.51 L1685.23 487.01 L1667.64 468.75 L1671.58 435.08 L1687 425.41 L1720.6801 445.89 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M561.24 794.95 L539.09 766.71 L508.48 772.43 L503.09 801.13 L515.12 813.83 L560.13 805.41 L561.24 794.95 Z"
      /><path d="M561.24 794.95 L539.09 766.71 L508.48 772.43 L503.09 801.13 L515.12 813.83 L560.13 805.41 L561.24 794.95 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M867.87 93.68 L861.92 111.23 L845.53 121.23 L841.19 120.69 L817.12 89.61 L817.93 78.12 L850.02 73.53 L867.87 93.68 Z"
      /><path d="M867.87 93.68 L861.92 111.23 L845.53 121.23 L841.19 120.69 L817.12 89.61 L817.93 78.12 L850.02 73.53 L867.87 93.68 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1812.2 175.39 L1825.73 176.97 L1843.1801 208.4 L1814.38 231.44 L1797.89 227.47 L1786.53 202.69 L1812.2 175.39 Z"
      /><path d="M1812.2 175.39 L1825.73 176.97 L1843.1801 208.4 L1814.38 231.44 L1797.89 227.47 L1786.53 202.69 L1812.2 175.39 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M352.34 59.64 L319.78 40.56 L292.32 56.26 L289.56 74.7 L309.03 99.61 L342.59 90.3 L352.34 59.64 Z"
      /><path d="M352.34 59.64 L319.78 40.56 L292.32 56.26 L289.56 74.7 L309.03 99.61 L342.59 90.3 L352.34 59.64 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M132.36 340.13 L129.93 366.74 L92.54 374.47 L80.6 363.28 L83.7 334.45 L111.6 323.27 L132.36 340.13 Z"
      /><path d="M132.36 340.13 L129.93 366.74 L92.54 374.47 L80.6 363.28 L83.7 334.45 L111.6 323.27 L132.36 340.13 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1301.5 413.86 L1256.78 379.3 L1246.5601 381.9 L1232.65 422.34 L1275.71 439.44 L1295.8101 428.11 L1301.76 415.95 L1301.5 413.86 Z"
      /><path d="M1301.5 413.86 L1256.78 379.3 L1246.5601 381.9 L1232.65 422.34 L1275.71 439.44 L1295.8101 428.11 L1301.76 415.95 L1301.5 413.86 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1027 245.77 L996.68 266.95 L996.58 282.81 L1014.29 297.03 L1040.0699 291.49 L1045.0601 257.25 L1027 245.77 Z"
      /><path d="M1027 245.77 L996.68 266.95 L996.58 282.81 L1014.29 297.03 L1040.0699 291.49 L1045.0601 257.25 L1027 245.77 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M63.76 161.34 L58.98 158.75 L37.2 164.54 L26.16 184.86 L40.69 205.45 L61.27 206.18 L72.29 195.66 L63.76 161.34 Z"
      /><path d="M63.76 161.34 L58.98 158.75 L37.2 164.54 L26.16 184.86 L40.69 205.45 L61.27 206.18 L72.29 195.66 L63.76 161.34 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1370.6801 333.49 L1342.34 320.92 L1330.4301 324.89 L1314.8 360.56 L1321.41 375.04 L1367.0601 382.52 L1370.6801 333.49 Z"
      /><path d="M1370.6801 333.49 L1342.34 320.92 L1330.4301 324.89 L1314.8 360.56 L1321.41 375.04 L1367.0601 382.52 L1370.6801 333.49 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M188.17 965.95 L144.08 932.08 L118.72 953.85 L156.38 1005.65 L182.37 991.96 L188.17 965.95 Z"
      /><path d="M188.17 965.95 L144.08 932.08 L118.72 953.85 L156.38 1005.65 L182.37 991.96 L188.17 965.95 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1793.23 652.88 L1777.33 678.61 L1746.17 679.46 L1738.15 671.08 L1747.77 631.46 L1773.97 629.96 L1793.23 652.88 Z"
      /><path d="M1793.23 652.88 L1777.33 678.61 L1746.17 679.46 L1738.15 671.08 L1747.77 631.46 L1773.97 629.96 L1793.23 652.88 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M772.12 71.31 L766.67 103.77 L790.8 115.41 L817.12 89.61 L817.93 78.12 L815.99 75.57 L772.12 71.31 Z"
      /><path d="M772.12 71.31 L766.67 103.77 L790.8 115.41 L817.12 89.61 L817.93 78.12 L815.99 75.57 L772.12 71.31 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M322.11 502.54 L362.19 522.77 L342.02 562.92 L306.5 552.95 L302.66 545.21 L312.66 508.28 L322.11 502.54 Z"
      /><path d="M322.11 502.54 L362.19 522.77 L342.02 562.92 L306.5 552.95 L302.66 545.21 L312.66 508.28 L322.11 502.54 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M99.28 476.33 L62.68 473.18 L48.21 496.29 L60.04 531.31 L81.57 536.16 L108.6 517.2 L99.28 476.33 Z"
      /><path d="M99.28 476.33 L62.68 473.18 L48.21 496.29 L60.04 531.31 L81.57 536.16 L108.6 517.2 L99.28 476.33 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1891.84 813.27 L1871.85 846.1 L1907.65 874.15 L1920 874.1 L1920 813.4 L1891.84 813.27 Z"
      /><path d="M1891.84 813.27 L1871.85 846.1 L1907.65 874.15 L1920 874.1 L1920 813.4 L1891.84 813.27 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1343.85 166.16 L1358.66 177.07 L1361.34 210.08 L1345.09 222.99 L1321.9 218.59 L1307.8199 181.41 L1312.6 172.23 L1343.85 166.16 Z"
      /><path d="M1343.85 166.16 L1358.66 177.07 L1361.34 210.08 L1345.09 222.99 L1321.9 218.59 L1307.8199 181.41 L1312.6 172.23 L1343.85 166.16 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M874.04 43.79 L891.85 60.73 L887.69 86.1 L867.87 93.68 L850.02 73.53 L861.76 43.84 L874.04 43.79 Z"
      /><path d="M874.04 43.79 L891.85 60.73 L887.69 86.1 L867.87 93.68 L850.02 73.53 L861.76 43.84 L874.04 43.79 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1584.79 54.22 L1584.61 79.64 L1578.48 86.3 L1537.76 88.95 L1529.3199 80.05 L1531.3101 51.27 L1550.34 39 L1584.79 54.22 Z"
      /><path d="M1584.79 54.22 L1584.61 79.64 L1578.48 86.3 L1537.76 88.95 L1529.3199 80.05 L1531.3101 51.27 L1550.34 39 L1584.79 54.22 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1498.1 173.88 L1529.48 194.77 L1531 214.44 L1502.23 223.75 L1481.5 201.87 L1492.88 174.36 L1498.1 173.88 Z"
      /><path d="M1498.1 173.88 L1529.48 194.77 L1531 214.44 L1502.23 223.75 L1481.5 201.87 L1492.88 174.36 L1498.1 173.88 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1389.28 691.76 L1408.5601 710.98 L1396.21 737.57 L1365.7 740.73 L1353.65 708.31 L1389.28 691.76 Z"
      /><path d="M1389.28 691.76 L1408.5601 710.98 L1396.21 737.57 L1365.7 740.73 L1353.65 708.31 L1389.28 691.76 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M581.12 475.22 L603.74 479.96 L608.37 528.57 L603.09 533.09 L576.22 530.26 L558.18 491.95 L581.12 475.22 Z"
      /><path d="M581.12 475.22 L603.74 479.96 L608.37 528.57 L603.09 533.09 L576.22 530.26 L558.18 491.95 L581.12 475.22 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M808.72 488.38 L789.56 498.82 L784.17 519.21 L815.8 545.16 L836.94 529.63 L835.42 501.16 L808.72 488.38 Z"
      /><path d="M808.72 488.38 L789.56 498.82 L784.17 519.21 L815.8 545.16 L836.94 529.63 L835.42 501.16 L808.72 488.38 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M395.27 299.37 L372.4 278.7 L342.87 298.13 L355.09 325.55 L391.92 313.05 L395.27 299.37 Z"
      /><path d="M395.27 299.37 L372.4 278.7 L342.87 298.13 L355.09 325.55 L391.92 313.05 L395.27 299.37 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1411.61 107.2 L1425.47 136.53 L1396.64 160.23 L1376.01 127.21 L1392.8101 103.68 L1411.61 107.2 Z"
      /><path d="M1411.61 107.2 L1425.47 136.53 L1396.64 160.23 L1376.01 127.21 L1392.8101 103.68 L1411.61 107.2 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M371.14 197.3 L405.09 215.07 L397.99 245.7 L372.4 256.04 L360.21 248.17 L356.34 208.67 L371.14 197.3 Z"
      /><path d="M371.14 197.3 L405.09 215.07 L397.99 245.7 L372.4 256.04 L360.21 248.17 L356.34 208.67 L371.14 197.3 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M615.33 981.56 L623.12 996.34 L610.14 1032.3101 L576.56 1028.41 L565.97 999.27 L568.12 993.83 L606.17 977.75 L615.33 981.56 Z"
      /><path d="M615.33 981.56 L623.12 996.34 L610.14 1032.3101 L576.56 1028.41 L565.97 999.27 L568.12 993.83 L606.17 977.75 L615.33 981.56 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M748.15 526.47 L764.23 530.54 L770.77 573.56 L746.56 582.18 L717.06 553.07 L748.15 526.47 Z"
      /><path d="M748.15 526.47 L764.23 530.54 L770.77 573.56 L746.56 582.18 L717.06 553.07 L748.15 526.47 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1170.48 994.51 L1194.54 1007.32 L1193.4 1033.36 L1165.22 1045.87 L1153.55 1038.74 L1147.26 1010.64 L1170.48 994.51 Z"
      /><path d="M1170.48 994.51 L1194.54 1007.32 L1193.4 1033.36 L1165.22 1045.87 L1153.55 1038.74 L1147.26 1010.64 L1170.48 994.51 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1732.9301 817.04 L1739.49 850.18 L1721.8101 869.43 L1694.48 865.57 L1682.53 844.74 L1694.37 815.1 L1712.6 808.1 L1732.9301 817.04 Z"
      /><path d="M1732.9301 817.04 L1739.49 850.18 L1721.8101 869.43 L1694.48 865.57 L1682.53 844.74 L1694.37 815.1 L1712.6 808.1 L1732.9301 817.04 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M50.45 77.12 L45.49 75.91 L24.94 91.28 L33.96 120.8 L55.06 124.7 L70.44 112.18 L50.45 77.12 Z"
      /><path d="M50.45 77.12 L45.49 75.91 L24.94 91.28 L33.96 120.8 L55.06 124.7 L70.44 112.18 L50.45 77.12 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1324.15 871.89 L1308.4399 878.52 L1300.1801 922.31 L1332.73 936.85 L1347.55 928.47 L1351.87 893.48 L1324.15 871.89 Z"
      /><path d="M1324.15 871.89 L1308.4399 878.52 L1300.1801 922.31 L1332.73 936.85 L1347.55 928.47 L1351.87 893.48 L1324.15 871.89 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M501.86 390.47 L497.9 399.91 L460.36 410.64 L442.7 373.13 L469.9 360.81 L501.86 390.47 Z"
      /><path d="M501.86 390.47 L497.9 399.91 L460.36 410.64 L442.7 373.13 L469.9 360.81 L501.86 390.47 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M724.19 306.84 L720.91 307.45 L701.55 336.31 L721.04 370.37 L738.98 372.29 L765.19 342.03 L764.33 336.19 L724.19 306.84 Z"
      /><path d="M724.19 306.84 L720.91 307.45 L701.55 336.31 L721.04 370.37 L738.98 372.29 L765.19 342.03 L764.33 336.19 L724.19 306.84 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1180.89 91.62 L1203.64 100.69 L1216.8 129.24 L1205.48 143.66 L1177.91 146.08 L1164.64 124.03 L1180.89 91.62 Z"
      /><path d="M1180.89 91.62 L1203.64 100.69 L1216.8 129.24 L1205.48 143.66 L1177.91 146.08 L1164.64 124.03 L1180.89 91.62 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M515.12 813.83 L503.09 801.13 L468.87 809.45 L465.8 839.93 L499.31 857.31 L514.29 851.73 L515.12 813.83 Z"
      /><path d="M515.12 813.83 L503.09 801.13 L468.87 809.45 L465.8 839.93 L499.31 857.31 L514.29 851.73 L515.12 813.83 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M576.56 1028.41 L610.14 1032.3101 L613.74 1037.5699 L606.3 1080 L572.9 1080 L565.94 1043 L576.56 1028.41 Z"
      /><path d="M576.56 1028.41 L610.14 1032.3101 L613.74 1037.5699 L606.3 1080 L572.9 1080 L565.94 1043 L576.56 1028.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1490.74 756.74 L1488.4 763.71 L1448.1899 780.85 L1433.46 760.75 L1445.65 737.03 L1476.84 732.65 L1490.74 756.74 Z"
      /><path d="M1490.74 756.74 L1488.4 763.71 L1448.1899 780.85 L1433.46 760.75 L1445.65 737.03 L1476.84 732.65 L1490.74 756.74 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1668.86 521.26 L1641.65 517.77 L1619.76 546.25 L1626.83 558.18 L1660.86 568.85 L1678.39 536.82 L1668.86 521.26 Z"
      /><path d="M1668.86 521.26 L1641.65 517.77 L1619.76 546.25 L1626.83 558.18 L1660.86 568.85 L1678.39 536.82 L1668.86 521.26 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1230.4 791.58 L1215.47 776.05 L1180.92 783.59 L1173.15 810.06 L1189.52 834.64 L1227.92 828.96 L1230.4 791.58 Z"
      /><path d="M1230.4 791.58 L1215.47 776.05 L1180.92 783.59 L1173.15 810.06 L1189.52 834.64 L1227.92 828.96 L1230.4 791.58 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M504.72 43.19 L513.88 50.08 L511.79 90.52 L481.54 99.1 L466.61 62.62 L473.44 48.47 L504.72 43.19 Z"
      /><path d="M504.72 43.19 L513.88 50.08 L511.79 90.52 L481.54 99.1 L466.61 62.62 L473.44 48.47 L504.72 43.19 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M103.2 624.55 L124.92 627.38 L143.06 665.78 L107.18 683.97 L79.12 653.1 L103.2 624.55 Z"
      /><path d="M103.2 624.55 L124.92 627.38 L143.06 665.78 L107.18 683.97 L79.12 653.1 L103.2 624.55 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1162.52 763.16 L1180.92 783.59 L1173.15 810.06 L1135.65 816.87 L1119.64 796.74 L1126.45 772.08 L1162.52 763.16 Z"
      /><path d="M1162.52 763.16 L1180.92 783.59 L1173.15 810.06 L1135.65 816.87 L1119.64 796.74 L1126.45 772.08 L1162.52 763.16 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M508.39 428.9 L536.26 437.55 L530.85 475.57 L500.61 477.86 L485.93 451.89 L508.39 428.9 Z"
      /><path d="M508.39 428.9 L536.26 437.55 L530.85 475.57 L500.61 477.86 L485.93 451.89 L508.39 428.9 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1247.62 610.72 L1217.8199 582.09 L1213.5 583.27 L1191.1899 614.86 L1205.76 641.62 L1236.6801 643.75 L1247.62 610.72 Z"
      /><path d="M1247.62 610.72 L1217.8199 582.09 L1213.5 583.27 L1191.1899 614.86 L1205.76 641.62 L1236.6801 643.75 L1247.62 610.72 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M845.53 121.23 L857.65 157.14 L828.67 171.16 L820.51 165.31 L815.87 138.01 L841.19 120.69 L845.53 121.23 Z"
      /><path d="M845.53 121.23 L857.65 157.14 L828.67 171.16 L820.51 165.31 L815.87 138.01 L841.19 120.69 L845.53 121.23 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M935.63 649.14 L917.29 648.78 L896.85 667.42 L899.97 695.86 L937.27 703.97 L949.66 684.81 L935.63 649.14 Z"
      /><path d="M935.63 649.14 L917.29 648.78 L896.85 667.42 L899.97 695.86 L937.27 703.97 L949.66 684.81 L935.63 649.14 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1122.3101 982.09 L1090.62 969.22 L1072.5601 985.78 L1076.9301 1005.25 L1107.39 1018.21 L1126.39 1002.39 L1122.3101 982.09 Z"
      /><path d="M1122.3101 982.09 L1090.62 969.22 L1072.5601 985.78 L1076.9301 1005.25 L1107.39 1018.21 L1126.39 1002.39 L1122.3101 982.09 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1875.39 1007.75 L1920 1015.5 L1920 1046.3 L1868.71 1046.59 L1859.1801 1024.62 L1875.39 1007.75 Z"
      /><path d="M1875.39 1007.75 L1920 1015.5 L1920 1046.3 L1868.71 1046.59 L1859.1801 1024.62 L1875.39 1007.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1279.84 969.78 L1312.23 983.15 L1307.52 1023.22 L1291.36 1029.33 L1258.26 1013.71 L1267.83 975.62 L1279.84 969.78 Z"
      /><path d="M1279.84 969.78 L1312.23 983.15 L1307.52 1023.22 L1291.36 1029.33 L1258.26 1013.71 L1267.83 975.62 L1279.84 969.78 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1300.3101 306.44 L1330.4301 324.89 L1314.8 360.56 L1276.92 352.59 L1269.7 324.31 L1300.3101 306.44 Z"
      /><path d="M1300.3101 306.44 L1330.4301 324.89 L1314.8 360.56 L1276.92 352.59 L1269.7 324.31 L1300.3101 306.44 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1285.3101 928.5 L1279.84 969.78 L1267.83 975.62 L1236.1801 961.05 L1236.63 931.17 L1262.11 918.05 L1285.3101 928.5 Z"
      /><path d="M1285.3101 928.5 L1279.84 969.78 L1267.83 975.62 L1236.1801 961.05 L1236.63 931.17 L1262.11 918.05 L1285.3101 928.5 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M274.19 494.38 L312.66 508.28 L302.66 545.21 L255.42 535.85 L250.79 526.44 L274.19 494.38 Z"
      /><path d="M274.19 494.38 L312.66 508.28 L302.66 545.21 L255.42 535.85 L250.79 526.44 L274.19 494.38 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1811.1801 1036.6 L1811 1080 L1753.5 1080 L1750.85 1025.92 L1776.91 1017.54 L1811.1801 1036.6 Z"
      /><path d="M1811.1801 1036.6 L1811 1080 L1753.5 1080 L1750.85 1025.92 L1776.91 1017.54 L1811.1801 1036.6 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M971.65 107.1 L969.87 62.79 L933.02 72.36 L930.11 83.67 L950.05 111.25 L971.65 107.1 Z"
      /><path d="M971.65 107.1 L969.87 62.79 L933.02 72.36 L930.11 83.67 L950.05 111.25 L971.65 107.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M804.87 660.08 L775.54 633.3 L766.62 634.9 L745.96 669.76 L773.1 694.79 L801.92 679.22 L804.87 660.08 Z"
      /><path d="M804.87 660.08 L775.54 633.3 L766.62 634.9 L745.96 669.76 L773.1 694.79 L801.92 679.22 L804.87 660.08 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1836.8199 836.81 L1790.5699 868.77 L1790.62 869.19 L1815.37 893.57 L1849.7 883.07 L1855.99 849.83 L1836.8199 836.81 Z"
      /><path d="M1836.8199 836.81 L1790.5699 868.77 L1790.62 869.19 L1815.37 893.57 L1849.7 883.07 L1855.99 849.83 L1836.8199 836.81 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1491.87 506.53 L1509.62 522.51 L1505.87 557.37 L1492.04 564.03 L1463.71 555.53 L1458.8101 525.16 L1491.87 506.53 Z"
      /><path d="M1491.87 506.53 L1509.62 522.51 L1505.87 557.37 L1492.04 564.03 L1463.71 555.53 L1458.8101 525.16 L1491.87 506.53 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1058.5 204.06 L1075.67 228.14 L1068.66 249.97 L1045.0601 257.25 L1027 245.77 L1022.59 227.53 L1034.9301 207.71 L1058.5 204.06 Z"
      /><path d="M1058.5 204.06 L1075.67 228.14 L1068.66 249.97 L1045.0601 257.25 L1027 245.77 L1022.59 227.53 L1034.9301 207.71 L1058.5 204.06 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1167.84 336.93 L1187.45 375.94 L1182.08 386.85 L1145 393.03 L1124.12 369.29 L1153.99 334.45 L1167.84 336.93 Z"
      /><path d="M1167.84 336.93 L1187.45 375.94 L1182.08 386.85 L1145 393.03 L1124.12 369.29 L1153.99 334.45 L1167.84 336.93 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1893.3 0 L1885.8199 31.69 L1857.29 35.44 L1852.85 30.64 L1853.9 0 L1893.3 0 Z"
      /><path d="M1893.3 0 L1885.8199 31.69 L1857.29 35.44 L1852.85 30.64 L1853.9 0 L1893.3 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1786.64 275.57 L1821.96 276.34 L1829.85 301.92 L1793.4399 323.28 L1774.54 302.74 L1786.64 275.57 Z"
      /><path d="M1786.64 275.57 L1821.96 276.34 L1829.85 301.92 L1793.4399 323.28 L1774.54 302.74 L1786.64 275.57 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M887.48 198.28 L875.55 191.79 L845.03 205.61 L854.45 240.71 L891.19 231.55 L887.48 198.28 Z"
      /><path d="M887.48 198.28 L875.55 191.79 L845.03 205.61 L854.45 240.71 L891.19 231.55 L887.48 198.28 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1441.92 139.24 L1425.47 136.53 L1396.64 160.23 L1396.53 160.83 L1412.03 185.89 L1438.21 188.04 L1454.28 158.16 L1441.92 139.24 Z"
      /><path d="M1441.92 139.24 L1425.47 136.53 L1396.64 160.23 L1396.53 160.83 L1412.03 185.89 L1438.21 188.04 L1454.28 158.16 L1441.92 139.24 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M29.07 914.03 L0 909.3 L0 971.9 L46.02 963.19 L51.16 949.59 L29.07 914.03 Z"
      /><path d="M29.07 914.03 L0 909.3 L0 971.9 L46.02 963.19 L51.16 949.59 L29.07 914.03 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M596.6 0 L550.9 0 L548.83 44.72 L558.26 52.58 L592.17 49.19 L599.97 40.53 L596.6 0 Z"
      /><path d="M596.6 0 L550.9 0 L548.83 44.72 L558.26 52.58 L592.17 49.19 L599.97 40.53 L596.6 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1873.03 615.44 L1920 619.5 L1920 652.9 L1872.83 657.57 L1863.5601 632.82 L1873.03 615.44 Z"
      /><path d="M1873.03 615.44 L1920 619.5 L1920 652.9 L1872.83 657.57 L1863.5601 632.82 L1873.03 615.44 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M942.13 273.59 L970.15 296.5 L966.56 319.17 L933.34 328.14 L919.47 307.06 L942.13 273.59 Z"
      /><path d="M942.13 273.59 L970.15 296.5 L966.56 319.17 L933.34 328.14 L919.47 307.06 L942.13 273.59 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M398.64 783.9 L364.81 789.89 L354.92 810.43 L367.78 832.42 L397.76 839.54 L411.99 829.27 L416.42 807.34 L398.64 783.9 Z"
      /><path d="M398.64 783.9 L364.81 789.89 L354.92 810.43 L367.78 832.42 L397.76 839.54 L411.99 829.27 L416.42 807.34 L398.64 783.9 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M545.94 491.11 L523.99 523.57 L546.29 553.73 L549.36 553.89 L576.22 530.26 L558.18 491.95 L545.94 491.11 Z"
      /><path d="M545.94 491.11 L523.99 523.57 L546.29 553.73 L549.36 553.89 L576.22 530.26 L558.18 491.95 L545.94 491.11 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1811.5 0 L1819.15 32.56 L1852.85 30.64 L1853.9 0 L1811.5 0 Z"
      /><path d="M1811.5 0 L1819.15 32.56 L1852.85 30.64 L1853.9 0 L1811.5 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M319.62 1049.8199 L320.2 1080 L256.6 1080 L256.47 1055.89 L282.63 1030.8199 L319.62 1049.8199 Z"
      /><path d="M319.62 1049.8199 L320.2 1080 L256.6 1080 L256.47 1055.89 L282.63 1030.8199 L319.62 1049.8199 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1776.02 461.75 L1757.36 485.75 L1769.09 511.96 L1804.05 508.7 L1815.5601 483.61 L1776.02 461.75 Z"
      /><path d="M1776.02 461.75 L1757.36 485.75 L1769.09 511.96 L1804.05 508.7 L1815.5601 483.61 L1776.02 461.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1774.55 37.37 L1787.1801 50.95 L1781.41 73.21 L1746.4 89.11 L1730.49 49.14 L1737.02 40.24 L1774.55 37.37 Z"
      /><path d="M1774.55 37.37 L1787.1801 50.95 L1781.41 73.21 L1746.4 89.11 L1730.49 49.14 L1737.02 40.24 L1774.55 37.37 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M951.33 501.24 L919.3 510.83 L919.85 546.25 L949.33 557.48 L971.5 529.71 L951.33 501.24 Z"
      /><path d="M951.33 501.24 L919.3 510.83 L919.85 546.25 L949.33 557.48 L971.5 529.71 L951.33 501.24 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M107.2 241.41 L92.69 281.25 L114.08 297.04 L139.51 285.26 L142.03 261.28 L107.2 241.41 Z"
      /><path d="M107.2 241.41 L92.69 281.25 L114.08 297.04 L139.51 285.26 L142.03 261.28 L107.2 241.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M463.98 1020.59 L481.43 1037.61 L477.8 1080 L432.6 1080 L429.65 1042 L457.29 1019.99 L463.98 1020.59 Z"
      /><path d="M463.98 1020.59 L481.43 1037.61 L477.8 1080 L432.6 1080 L429.65 1042 L457.29 1019.99 L463.98 1020.59 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M549.6 393.46 L553.34 428.25 L536.26 437.55 L508.39 428.9 L497.9 399.91 L501.86 390.47 L516.64 381.26 L549.6 393.46 Z"
      /><path d="M549.6 393.46 L553.34 428.25 L536.26 437.55 L508.39 428.9 L497.9 399.91 L501.86 390.47 L516.64 381.26 L549.6 393.46 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M906.46 596.44 L938.43 597.59 L951.84 632.89 L935.63 649.14 L917.29 648.78 L894.75 610.04 L906.46 596.44 Z"
      /><path d="M906.46 596.44 L938.43 597.59 L951.84 632.89 L935.63 649.14 L917.29 648.78 L894.75 610.04 L906.46 596.44 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M508.39 428.9 L497.9 399.91 L460.36 410.64 L453.87 424.48 L468.84 449.46 L485.93 451.89 L508.39 428.9 Z"
      /><path d="M508.39 428.9 L497.9 399.91 L460.36 410.64 L453.87 424.48 L468.84 449.46 L485.93 451.89 L508.39 428.9 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1842.27 962.59 L1825.72 978.93 L1836.99 1019.63 L1859.1801 1024.62 L1875.39 1007.75 L1876.58 972.05 L1875.54 970.71 L1842.27 962.59 Z"
      /><path d="M1842.27 962.59 L1825.72 978.93 L1836.99 1019.63 L1859.1801 1024.62 L1875.39 1007.75 L1876.58 972.05 L1875.54 970.71 L1842.27 962.59 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M209.89 216.96 L180.14 196.88 L154.2 216.22 L162.79 246.69 L175.47 250.2 L209.08 220.61 L209.89 216.96 Z"
      /><path d="M209.89 216.96 L180.14 196.88 L154.2 216.22 L162.79 246.69 L175.47 250.2 L209.08 220.61 L209.89 216.96 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M174.56 430.14 L160.69 427.88 L125.38 460.08 L165.34 493.73 L173.17 487.85 L183.79 442.98 L174.56 430.14 Z"
      /><path d="M174.56 430.14 L160.69 427.88 L125.38 460.08 L165.34 493.73 L173.17 487.85 L183.79 442.98 L174.56 430.14 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1256.1 0 L1293.8 0 L1298.71 36.45 L1285.28 51.19 L1255.8 43.42 L1256.1 0 Z"
      /><path d="M1256.1 0 L1293.8 0 L1298.71 36.45 L1285.28 51.19 L1255.8 43.42 L1256.1 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1448 687.18 L1483.0601 713.66 L1476.84 732.65 L1445.65 737.03 L1428.8 708.05 L1443.29 688.24 L1448 687.18 Z"
      /><path d="M1448 687.18 L1483.0601 713.66 L1476.84 732.65 L1445.65 737.03 L1428.8 708.05 L1443.29 688.24 L1448 687.18 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M92.46 196.84 L72.29 195.66 L61.27 206.18 L69.76 236.99 L106.32 239.18 L109.45 229.29 L92.46 196.84 Z"
      /><path d="M92.46 196.84 L72.29 195.66 L61.27 206.18 L69.76 236.99 L106.32 239.18 L109.45 229.29 L92.46 196.84 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M847.69 697.79 L883.61 711.9 L885.39 735.96 L859.86 756.17 L840.97 752.41 L826.4 722.82 L832.16 705.26 L847.69 697.79 Z"
      /><path d="M847.69 697.79 L883.61 711.9 L885.39 735.96 L859.86 756.17 L840.97 752.41 L826.4 722.82 L832.16 705.26 L847.69 697.79 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1920 753.5 L1920 813.4 L1891.84 813.27 L1871.04 788.85 L1898.05 754.18 L1920 753.5 Z"
      /><path d="M1920 753.5 L1920 813.4 L1891.84 813.27 L1871.04 788.85 L1898.05 754.18 L1920 753.5 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1458.8101 525.16 L1438.78 514.74 L1404.45 537.68 L1403.91 540.07 L1418.89 564.96 L1446.77 570.84 L1463.71 555.53 L1458.8101 525.16 Z"
      /><path d="M1458.8101 525.16 L1438.78 514.74 L1404.45 537.68 L1403.91 540.07 L1418.89 564.96 L1446.77 570.84 L1463.71 555.53 L1458.8101 525.16 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M847.78 361.89 L819.16 351.79 L799.89 362.43 L795.81 396.68 L831.79 409.55 L852.23 396.25 L847.78 361.89 Z"
      /><path d="M847.78 361.89 L819.16 351.79 L799.89 362.43 L795.81 396.68 L831.79 409.55 L852.23 396.25 L847.78 361.89 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1172.9 230.44 L1219.04 239.61 L1213.51 275.7 L1192.9301 287.35 L1173.45 277.16 L1166.47 240.71 L1172.9 230.44 Z"
      /><path d="M1172.9 230.44 L1219.04 239.61 L1213.51 275.7 L1192.9301 287.35 L1173.45 277.16 L1166.47 240.71 L1172.9 230.44 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M831.41 444.97 L811.74 455.03 L808.72 488.38 L835.42 501.16 L858.21 485.7 L856.62 456.72 L831.41 444.97 Z"
      /><path d="M831.41 444.97 L811.74 455.03 L808.72 488.38 L835.42 501.16 L858.21 485.7 L856.62 456.72 L831.41 444.97 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M775.3 981.35 L766.93 949.45 L727.4 954.25 L717.95 983.19 L752.37 1001.03 L775.3 981.35 Z"
      /><path d="M775.3 981.35 L766.93 949.45 L727.4 954.25 L717.95 983.19 L752.37 1001.03 L775.3 981.35 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1192.9301 287.35 L1173.45 277.16 L1139.72 294.11 L1136.0699 308.24 L1153.99 334.45 L1167.84 336.93 L1194.4301 316.57 L1192.9301 287.35 Z"
      /><path d="M1192.9301 287.35 L1173.45 277.16 L1139.72 294.11 L1136.0699 308.24 L1153.99 334.45 L1167.84 336.93 L1194.4301 316.57 L1192.9301 287.35 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1660.86 568.85 L1662.66 573.54 L1644.1801 608.46 L1613.64 596.12 L1626.83 558.18 L1660.86 568.85 Z"
      /><path d="M1660.86 568.85 L1662.66 573.54 L1644.1801 608.46 L1613.64 596.12 L1626.83 558.18 L1660.86 568.85 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M271.25 944.86 L302.93 965.68 L301.79 990.77 L281.63 1007.9 L246.3 991.33 L244.09 968.82 L271.25 944.86 Z"
      /><path d="M271.25 944.86 L302.93 965.68 L301.79 990.77 L281.63 1007.9 L246.3 991.33 L244.09 968.82 L271.25 944.86 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1442.97 84.35 L1458.88 114.22 L1441.92 139.24 L1425.47 136.53 L1411.61 107.2 L1439.85 83.03 L1442.97 84.35 Z"
      /><path d="M1442.97 84.35 L1458.88 114.22 L1441.92 139.24 L1425.47 136.53 L1411.61 107.2 L1439.85 83.03 L1442.97 84.35 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M427.02 701.99 L446.42 718.75 L439.41 752.39 L407.52 758.11 L390.45 735.12 L401.54 708.16 L427.02 701.99 Z"
      /><path d="M427.02 701.99 L446.42 718.75 L439.41 752.39 L407.52 758.11 L390.45 735.12 L401.54 708.16 L427.02 701.99 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1787.78 596.18 L1773.97 629.96 L1747.77 631.46 L1736.39 621.14 L1743.5699 581.99 L1748.92 579.08 L1787.78 596.18 Z"
      /><path d="M1787.78 596.18 L1773.97 629.96 L1747.77 631.46 L1736.39 621.14 L1743.5699 581.99 L1748.92 579.08 L1787.78 596.18 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1242.08 509.3 L1263.67 525.19 L1258.97 556.57 L1229.52 563.84 L1213.3199 523.34 L1242.08 509.3 Z"
      /><path d="M1242.08 509.3 L1263.67 525.19 L1258.97 556.57 L1229.52 563.84 L1213.3199 523.34 L1242.08 509.3 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1552.85 991.24 L1522.3 971.41 L1491.51 980.97 L1482.92 999.72 L1488.02 1020.63 L1520.9301 1038.36 L1552.96 1018.15 L1557.6 1005.65 L1552.85 991.24 Z"
      /><path d="M1552.85 991.24 L1522.3 971.41 L1491.51 980.97 L1482.92 999.72 L1488.02 1020.63 L1520.9301 1038.36 L1552.96 1018.15 L1557.6 1005.65 L1552.85 991.24 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1332.73 936.85 L1300.1801 922.31 L1285.3101 928.5 L1279.84 969.78 L1312.23 983.15 L1328.4 974.22 L1332.73 936.85 Z"
      /><path d="M1332.73 936.85 L1300.1801 922.31 L1285.3101 928.5 L1279.84 969.78 L1312.23 983.15 L1328.4 974.22 L1332.73 936.85 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1680.03 345.36 L1656.22 320.97 L1624.0601 329.35 L1619 339.09 L1639.16 379.22 L1664.0699 374.41 L1680.03 345.36 Z"
      /><path d="M1680.03 345.36 L1656.22 320.97 L1624.0601 329.35 L1619 339.09 L1639.16 379.22 L1664.0699 374.41 L1680.03 345.36 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M305.94 656.28 L277.53 626.61 L260.22 632.73 L254.08 670.77 L289.8 681.11 L305.94 656.28 Z"
      /><path d="M305.94 656.28 L277.53 626.61 L260.22 632.73 L254.08 670.77 L289.8 681.11 L305.94 656.28 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1359.45 428.61 L1353.6801 457.3 L1325.74 474.37 L1323.37 473.87 L1295.8101 428.11 L1301.76 415.95 L1359.45 428.61 Z"
      /><path d="M1359.45 428.61 L1353.6801 457.3 L1325.74 474.37 L1323.37 473.87 L1295.8101 428.11 L1301.76 415.95 L1359.45 428.61 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1573.34 437.05 L1525.45 417.45 L1512.49 423.55 L1519.9399 468.17 L1547.08 479.64 L1565.23 469.67 L1573.34 437.05 Z"
      /><path d="M1573.34 437.05 L1525.45 417.45 L1512.49 423.55 L1519.9399 468.17 L1547.08 479.64 L1565.23 469.67 L1573.34 437.05 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1415.4399 656.69 L1443.29 688.24 L1428.8 708.05 L1408.5601 710.98 L1389.28 691.76 L1391.21 661.61 L1415.4399 656.69 Z"
      /><path d="M1415.4399 656.69 L1443.29 688.24 L1428.8 708.05 L1408.5601 710.98 L1389.28 691.76 L1391.21 661.61 L1415.4399 656.69 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M24.94 91.28 L0 88 L0 138.6 L13.63 138.41 L33.96 120.8 L24.94 91.28 Z"
      /><path d="M24.94 91.28 L0 88 L0 138.6 L13.63 138.41 L33.96 120.8 L24.94 91.28 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1446.77 570.84 L1451.4 597.09 L1428.64 619.02 L1398.9399 601.52 L1418.89 564.96 L1446.77 570.84 Z"
      /><path d="M1446.77 570.84 L1451.4 597.09 L1428.64 619.02 L1398.9399 601.52 L1418.89 564.96 L1446.77 570.84 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M679.28 653.48 L661.97 640.38 L640.93 644.84 L627.19 672.96 L643.45 697.68 L667.74 699.74 L677.35 691.73 L679.28 653.48 Z"
      /><path d="M679.28 653.48 L661.97 640.38 L640.93 644.84 L627.19 672.96 L643.45 697.68 L667.74 699.74 L677.35 691.73 L679.28 653.48 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1620.46 151.82 L1657.4399 153.61 L1665.4 187.98 L1645.08 198.8 L1617.89 189.49 L1611.35 170.9 L1620.46 151.82 Z"
      /><path d="M1620.46 151.82 L1657.4399 153.61 L1665.4 187.98 L1645.08 198.8 L1617.89 189.49 L1611.35 170.9 L1620.46 151.82 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M543.75 336.54 L551.09 337.73 L575.42 369.03 L575.53 370.92 L549.6 393.46 L516.64 381.26 L520.45 351.88 L543.75 336.54 Z"
      /><path d="M543.75 336.54 L551.09 337.73 L575.42 369.03 L575.53 370.92 L549.6 393.46 L516.64 381.26 L520.45 351.88 L543.75 336.54 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M820.14 307.27 L806.07 297.96 L790.1 300.51 L764.33 336.19 L765.19 342.03 L799.89 362.43 L819.16 351.79 L820.14 307.27 Z"
      /><path d="M820.14 307.27 L806.07 297.96 L790.1 300.51 L764.33 336.19 L765.19 342.03 L799.89 362.43 L819.16 351.79 L820.14 307.27 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M360.13 389.86 L362.87 413.88 L335.43 429.57 L311.67 414.39 L312.2 390.58 L335.6 377 L360.13 389.86 Z"
      /><path d="M360.13 389.86 L362.87 413.88 L335.43 429.57 L311.67 414.39 L312.2 390.58 L335.6 377 L360.13 389.86 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M583.07 897.17 L574.09 878.67 L538.17 883.31 L529.74 907.42 L566.49 927.27 L583.07 897.17 Z"
      /><path d="M583.07 897.17 L574.09 878.67 L538.17 883.31 L529.74 907.42 L566.49 927.27 L583.07 897.17 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1274.58 833.23 L1280.14 867.75 L1257.53 882.86 L1233.39 874.91 L1230.13 831.05 L1274.58 833.23 Z"
      /><path d="M1274.58 833.23 L1280.14 867.75 L1257.53 882.86 L1233.39 874.91 L1230.13 831.05 L1274.58 833.23 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M182.37 991.96 L219.29 1017.45 L219.85 1026.79 L183.08 1066.5601 L150.41 1017.44 L156.38 1005.65 L182.37 991.96 Z"
      /><path d="M182.37 991.96 L219.29 1017.45 L219.85 1026.79 L183.08 1066.5601 L150.41 1017.44 L156.38 1005.65 L182.37 991.96 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1420.36 1008.66 L1420.17 1024.54 L1390.3199 1049.8101 L1357.4 1026.0601 L1365.36 991.44 L1372.8199 987.48 L1420.36 1008.66 Z"
      /><path d="M1420.36 1008.66 L1420.17 1024.54 L1390.3199 1049.8101 L1357.4 1026.0601 L1365.36 991.44 L1372.8199 987.48 L1420.36 1008.66 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1829.85 301.92 L1839.52 307.88 L1844.87 345.48 L1815.33 354.62 L1793.33 339.37 L1793.4399 323.28 L1829.85 301.92 Z"
      /><path d="M1829.85 301.92 L1839.52 307.88 L1844.87 345.48 L1815.33 354.62 L1793.33 339.37 L1793.4399 323.28 L1829.85 301.92 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M253.71 770.18 L284.77 801.54 L267.97 830.51 L230.73 824.75 L232.91 786.42 L253.71 770.18 Z"
      /><path d="M253.71 770.18 L284.77 801.54 L267.97 830.51 L230.73 824.75 L232.91 786.42 L253.71 770.18 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M770.7 0 L743.3 0 L738.99 52.64 L764.15 58.04 L781.96 35.92 L770.7 0 Z"
      /><path d="M770.7 0 L743.3 0 L738.99 52.64 L764.15 58.04 L781.96 35.92 L770.7 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1013.07 76.53 L1014.8 87.25 L989.56 116.82 L971.65 107.1 L969.87 62.79 L975.05 56.27 L982.91 54.64 L1013.07 76.53 Z"
      /><path d="M1013.07 76.53 L1014.8 87.25 L989.56 116.82 L971.65 107.1 L969.87 62.79 L975.05 56.27 L982.91 54.64 L1013.07 76.53 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1046.26 723.17 L1074 756.27 L1066.3 774.35 L1032.83 779.36 L1014.68 747.47 L1046.26 723.17 Z"
      /><path d="M1046.26 723.17 L1074 756.27 L1066.3 774.35 L1032.83 779.36 L1014.68 747.47 L1046.26 723.17 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1328.4 974.22 L1312.23 983.15 L1307.52 1023.22 L1333.4 1037.48 L1357.4 1026.0601 L1365.36 991.44 L1328.4 974.22 Z"
      /><path d="M1328.4 974.22 L1312.23 983.15 L1307.52 1023.22 L1333.4 1037.48 L1357.4 1026.0601 L1365.36 991.44 L1328.4 974.22 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1106.1 96.92 L1125.02 103.95 L1134.52 122.63 L1122.88 147.29 L1092.24 149.06 L1081.42 130.1 L1091.0601 103.39 L1106.1 96.92 Z"
      /><path d="M1106.1 96.92 L1125.02 103.95 L1134.52 122.63 L1122.88 147.29 L1092.24 149.06 L1081.42 130.1 L1091.0601 103.39 L1106.1 96.92 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M619.77 429.11 L603.61 419.04 L571.04 434.9 L581.12 475.22 L603.74 479.96 L621.16 470.64 L619.77 429.11 Z"
      /><path d="M619.77 429.11 L603.61 419.04 L571.04 434.9 L581.12 475.22 L603.74 479.96 L621.16 470.64 L619.77 429.11 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M428.61 101.91 L424.42 105.93 L439.04 147.17 L479.43 132.99 L478.6 103.61 L428.61 101.91 Z"
      /><path d="M428.61 101.91 L424.42 105.93 L439.04 147.17 L479.43 132.99 L478.6 103.61 L428.61 101.91 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1757.36 485.75 L1769.09 511.96 L1758.04 536.89 L1721.35 529.12 L1716.37 485.51 L1719.91 482.23 L1757.36 485.75 Z"
      /><path d="M1757.36 485.75 L1769.09 511.96 L1758.04 536.89 L1721.35 529.12 L1716.37 485.51 L1719.91 482.23 L1757.36 485.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M592.11 770.57 L617.67 783.67 L616.16 816.42 L610.85 821.19 L564.3 812.76 L560.13 805.41 L561.24 794.95 L592.11 770.57 Z"
      /><path d="M592.11 770.57 L617.67 783.67 L616.16 816.42 L610.85 821.19 L564.3 812.76 L560.13 805.41 L561.24 794.95 L592.11 770.57 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M985.61 219.15 L939.82 209.71 L939.74 209.75 L936.75 217.86 L951.94 254.88 L977.87 248.46 L985.66 219.24 L985.61 219.15 Z"
      /><path d="M985.61 219.15 L939.82 209.71 L939.74 209.75 L936.75 217.86 L951.94 254.88 L977.87 248.46 L985.66 219.24 L985.61 219.15 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1779.5 0 L1774.55 37.37 L1787.1801 50.95 L1811.0699 45.68 L1819.15 32.56 L1811.5 0 L1779.5 0 Z"
      /><path d="M1779.5 0 L1774.55 37.37 L1787.1801 50.95 L1811.0699 45.68 L1819.15 32.56 L1811.5 0 L1779.5 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M61.27 206.18 L69.76 236.99 L56.14 252.55 L44.7 253.81 L25.48 227.98 L40.69 205.45 L61.27 206.18 Z"
      /><path d="M61.27 206.18 L69.76 236.99 L56.14 252.55 L44.7 253.81 L25.48 227.98 L40.69 205.45 L61.27 206.18 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1349.85 82.34 L1340.75 119.08 L1317.6899 119.5 L1295.78 83.87 L1339.8101 69.47 L1349.85 82.34 Z"
      /><path d="M1349.85 82.34 L1340.75 119.08 L1317.6899 119.5 L1295.78 83.87 L1339.8101 69.47 L1349.85 82.34 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1170.8 215.28 L1172.9 230.44 L1166.47 240.71 L1125.11 246.75 L1111.26 219.53 L1117.75 201.94 L1127.17 196.34 L1170.8 215.28 Z"
      /><path d="M1170.8 215.28 L1172.9 230.44 L1166.47 240.71 L1125.11 246.75 L1111.26 219.53 L1117.75 201.94 L1127.17 196.34 L1170.8 215.28 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1748.77 351.56 L1740.16 313.65 L1710.03 315.54 L1693.98 342.71 L1722.5699 367.48 L1748.77 351.56 Z"
      /><path d="M1748.77 351.56 L1740.16 313.65 L1710.03 315.54 L1693.98 342.71 L1722.5699 367.48 L1748.77 351.56 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M317.91 294.11 L287.48 275.3 L278.6 277.5 L262.07 313.98 L263.24 316.12 L301.57 327.21 L317.91 294.11 Z"
      /><path d="M317.91 294.11 L287.48 275.3 L278.6 277.5 L262.07 313.98 L263.24 316.12 L301.57 327.21 L317.91 294.11 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1246.76 290.96 L1213.51 275.7 L1192.9301 287.35 L1194.4301 316.57 L1223.54 331.81 L1250.73 314.49 L1246.76 290.96 Z"
      /><path d="M1246.76 290.96 L1213.51 275.7 L1192.9301 287.35 L1194.4301 316.57 L1223.54 331.81 L1250.73 314.49 L1246.76 290.96 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M707.76 211.4 L704.5 242.05 L689.93 254.6 L644.06 234.27 L642.48 212.11 L673.51 192.33 L707.76 211.4 Z"
      /><path d="M707.76 211.4 L704.5 242.05 L689.93 254.6 L644.06 234.27 L642.48 212.11 L673.51 192.33 L707.76 211.4 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1432.4 994.24 L1482.92 999.72 L1488.02 1020.63 L1455.34 1052.53 L1420.17 1024.54 L1420.36 1008.66 L1432.4 994.24 Z"
      /><path d="M1432.4 994.24 L1482.92 999.72 L1488.02 1020.63 L1455.34 1052.53 L1420.17 1024.54 L1420.36 1008.66 L1432.4 994.24 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1830.84 815.43 L1836.8199 836.81 L1790.5699 868.77 L1780.6801 856.76 L1785.6899 810.85 L1801.16 803.13 L1830.84 815.43 Z"
      /><path d="M1830.84 815.43 L1836.8199 836.81 L1790.5699 868.77 L1780.6801 856.76 L1785.6899 810.85 L1801.16 803.13 L1830.84 815.43 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1463.71 555.53 L1446.77 570.84 L1451.4 597.09 L1488.24 611.46 L1492.04 564.03 L1463.71 555.53 Z"
      /><path d="M1463.71 555.53 L1446.77 570.84 L1451.4 597.09 L1488.24 611.46 L1492.04 564.03 L1463.71 555.53 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M371.18 519.93 L397.2 546.84 L393.92 579.01 L388.46 584.77 L347.82 574.24 L342.02 562.92 L362.19 522.77 L371.18 519.93 Z"
      /><path d="M371.18 519.93 L397.2 546.84 L393.92 579.01 L388.46 584.77 L347.82 574.24 L342.02 562.92 L362.19 522.77 L371.18 519.93 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1825.72 978.93 L1836.99 1019.63 L1811.1801 1036.6 L1776.91 1017.54 L1792.24 976.03 L1825.72 978.93 Z"
      /><path d="M1825.72 978.93 L1836.99 1019.63 L1811.1801 1036.6 L1776.91 1017.54 L1792.24 976.03 L1825.72 978.93 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1871.54 905.64 L1849.7 883.07 L1815.37 893.57 L1814.84 921.49 L1837.64 936.51 L1871.77 911.85 L1871.54 905.64 Z"
      /><path d="M1871.54 905.64 L1849.7 883.07 L1815.37 893.57 L1814.84 921.49 L1837.64 936.51 L1871.77 911.85 L1871.54 905.64 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1310.14 750.49 L1325.1801 761.94 L1327 792.95 L1305.04 814.21 L1289.9 814.35 L1270.35 783.27 L1277.4301 760.51 L1310.14 750.49 Z"
      /><path d="M1310.14 750.49 L1325.1801 761.94 L1327 792.95 L1305.04 814.21 L1289.9 814.35 L1270.35 783.27 L1277.4301 760.51 L1310.14 750.49 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M77 0 L32.9 0 L39.5 36.03 L73.08 32.67 L77 0 Z"
      /><path d="M77 0 L32.9 0 L39.5 36.03 L73.08 32.67 L77 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M989 857.11 L1004.14 863.84 L1010.04 907.21 L1003.63 913.93 L971 913.61 L954.76 881.86 L989 857.11 Z"
      /><path d="M989 857.11 L1004.14 863.84 L1010.04 907.21 L1003.63 913.93 L971 913.61 L954.76 881.86 L989 857.11 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1650.98 275.8 L1665.37 291.54 L1656.22 320.97 L1624.0601 329.35 L1607.84 291.38 L1610.75 284.8 L1650.98 275.8 Z"
      /><path d="M1650.98 275.8 L1665.37 291.54 L1656.22 320.97 L1624.0601 329.35 L1607.84 291.38 L1610.75 284.8 L1650.98 275.8 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1721.35 529.12 L1716.37 485.51 L1685.23 487.01 L1668.86 521.26 L1678.39 536.82 L1706.4301 541.91 L1721.35 529.12 Z"
      /><path d="M1721.35 529.12 L1716.37 485.51 L1685.23 487.01 L1668.86 521.26 L1678.39 536.82 L1706.4301 541.91 L1721.35 529.12 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1694.49 696.82 L1674.28 687.65 L1647.64 702.72 L1650.48 725.5 L1669.97 735.46 L1699.78 713.58 L1694.49 696.82 Z"
      /><path d="M1694.49 696.82 L1674.28 687.65 L1647.64 702.72 L1650.48 725.5 L1669.97 735.46 L1699.78 713.58 L1694.49 696.82 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1005.05 483.78 L966.19 472.72 L960.92 475.28 L951.33 501.24 L971.5 529.71 L989.06 530.77 L1015.37 504.89 L1005.05 483.78 Z"
      /><path d="M1005.05 483.78 L966.19 472.72 L960.92 475.28 L951.33 501.24 L971.5 529.71 L989.06 530.77 L1015.37 504.89 L1005.05 483.78 Z" style="fill:rgb(0,225,0); stroke:none;"
      /><path style="fill:none;" d="M910.29 455.31 L899.95 498.36 L887.61 501.45 L858.21 485.7 L856.62 456.72 L880.43 441.82 L910.29 455.31 Z"
      /><path d="M910.29 455.31 L899.95 498.36 L887.61 501.45 L858.21 485.7 L856.62 456.72 L880.43 441.82 L910.29 455.31 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1019.72 803.99 L998.67 805.52 L980.08 830.88 L989 857.11 L1004.14 863.84 L1033.1801 852.13 L1038.8 827.94 L1019.72 803.99 Z"
      /><path d="M1019.72 803.99 L998.67 805.52 L980.08 830.88 L989 857.11 L1004.14 863.84 L1033.1801 852.13 L1038.8 827.94 L1019.72 803.99 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1879.78 73.59 L1855.91 61.41 L1834.02 74.78 L1830.99 86.85 L1865.0699 111.69 L1883.78 92.87 L1879.78 73.59 Z"
      /><path d="M1879.78 73.59 L1855.91 61.41 L1834.02 74.78 L1830.99 86.85 L1865.0699 111.69 L1883.78 92.87 L1879.78 73.59 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1382.79 83.73 L1392.8101 103.68 L1376.01 127.21 L1349.73 128.01 L1340.75 119.08 L1349.85 82.34 L1382.79 83.73 Z"
      /><path d="M1382.79 83.73 L1392.8101 103.68 L1376.01 127.21 L1349.73 128.01 L1340.75 119.08 L1349.85 82.34 L1382.79 83.73 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M266.9 0 L210 0 L209.56 30.24 L231.98 51.27 L265.18 32.15 L266.9 0 Z"
      /><path d="M266.9 0 L210 0 L209.56 30.24 L231.98 51.27 L265.18 32.15 L266.9 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1735.35 904.98 L1756.72 909.05 L1777.9301 942.05 L1775.95 952.44 L1725.75 972.5 L1709.85 928.62 L1735.35 904.98 Z"
      /><path d="M1735.35 904.98 L1756.72 909.05 L1777.9301 942.05 L1775.95 952.44 L1725.75 972.5 L1709.85 928.62 L1735.35 904.98 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M773.1 694.79 L745.96 669.76 L732.37 671.54 L715.15 697.93 L724.43 726.1 L733.93 731.16 L770.25 716.02 L773.1 694.79 Z"
      /><path d="M773.1 694.79 L745.96 669.76 L732.37 671.54 L715.15 697.93 L724.43 726.1 L733.93 731.16 L770.25 716.02 L773.1 694.79 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1413.1801 760.19 L1389.11 792.48 L1380.71 792.56 L1359.77 751.15 L1365.7 740.73 L1396.21 737.57 L1413.1801 760.19 Z"
      /><path d="M1413.1801 760.19 L1389.11 792.48 L1380.71 792.56 L1359.77 751.15 L1365.7 740.73 L1396.21 737.57 L1413.1801 760.19 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1674.46 131.47 L1657.4399 153.61 L1665.4 187.98 L1677.91 193.05 L1707.4 184.11 L1710.73 178.37 L1704.8199 146.48 L1674.46 131.47 Z"
      /><path d="M1674.46 131.47 L1657.4399 153.61 L1665.4 187.98 L1677.91 193.05 L1707.4 184.11 L1710.73 178.37 L1704.8199 146.48 L1674.46 131.47 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M219.85 1026.79 L256.47 1055.89 L256.6 1080 L181.8 1080 L183.08 1066.5601 L219.85 1026.79 Z"
      /><path d="M219.85 1026.79 L256.47 1055.89 L256.6 1080 L181.8 1080 L183.08 1066.5601 L219.85 1026.79 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M704.5 242.05 L752.48 261.1 L752.9 269.91 L724.19 306.84 L720.91 307.45 L687.27 278.18 L689.93 254.6 L704.5 242.05 Z"
      /><path d="M704.5 242.05 L752.48 261.1 L752.9 269.91 L724.19 306.84 L720.91 307.45 L687.27 278.18 L689.93 254.6 L704.5 242.05 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M145.37 759.14 L183.51 774.17 L178 810.2 L144.38 830.79 L123.38 815.88 L120.99 777.28 L145.37 759.14 Z"
      /><path d="M145.37 759.14 L183.51 774.17 L178 810.2 L144.38 830.79 L123.38 815.88 L120.99 777.28 L145.37 759.14 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M760.31 156.27 L771.29 159.63 L782.12 175.02 L781.08 195.16 L758.09 212.02 L726.75 198.67 L729.47 170.58 L760.31 156.27 Z"
      /><path d="M760.31 156.27 L771.29 159.63 L782.12 175.02 L781.08 195.16 L758.09 212.02 L726.75 198.67 L729.47 170.58 L760.31 156.27 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M917.29 648.78 L894.75 610.04 L879.82 612.59 L858.82 652.73 L896.85 667.42 L917.29 648.78 Z"
      /><path d="M917.29 648.78 L894.75 610.04 L879.82 612.59 L858.82 652.73 L896.85 667.42 L917.29 648.78 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M852.23 396.25 L877.75 406.2 L880.43 441.82 L856.62 456.72 L831.41 444.97 L831.79 409.55 L852.23 396.25 Z"
      /><path d="M852.23 396.25 L877.75 406.2 L880.43 441.82 L856.62 456.72 L831.41 444.97 L831.79 409.55 L852.23 396.25 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1054.03 393.2 L1023.33 392.45 L1009.14 429.87 L1024 447.36 L1049.77 448.68 L1066.8199 406.2 L1054.03 393.2 Z"
      /><path d="M1054.03 393.2 L1023.33 392.45 L1009.14 429.87 L1024 447.36 L1049.77 448.68 L1066.8199 406.2 L1054.03 393.2 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M920.81 399.33 L899.98 393.03 L877.75 406.2 L880.43 441.82 L910.29 455.31 L921.15 450.84 L933.12 420.38 L920.81 399.33 Z"
      /><path d="M920.81 399.33 L899.98 393.03 L877.75 406.2 L880.43 441.82 L910.29 455.31 L921.15 450.84 L933.12 420.38 L920.81 399.33 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M405.74 337.96 L391.92 313.05 L355.09 325.55 L351.99 336.07 L385.1 362.8 L405.74 337.96 Z"
      /><path d="M405.74 337.96 L391.92 313.05 L355.09 325.55 L351.99 336.07 L385.1 362.8 L405.74 337.96 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M13.63 138.41 L37.2 164.54 L26.16 184.86 L0 186.2 L0 138.6 L13.63 138.41 Z"
      /><path d="M13.63 138.41 L37.2 164.54 L26.16 184.86 L0 186.2 L0 138.6 L13.63 138.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M698.66 781.84 L714.19 786.36 L726.71 813.38 L708.1 839.98 L666.53 822.38 L671.18 799.59 L698.66 781.84 Z"
      /><path d="M698.66 781.84 L714.19 786.36 L726.71 813.38 L708.1 839.98 L666.53 822.38 L671.18 799.59 L698.66 781.84 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1815.37 893.57 L1790.62 869.19 L1756.72 909.05 L1777.9301 942.05 L1814.84 921.49 L1815.37 893.57 Z"
      /><path d="M1815.37 893.57 L1790.62 869.19 L1756.72 909.05 L1777.9301 942.05 L1814.84 921.49 L1815.37 893.57 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M807.25 836.89 L828.26 866.42 L810.8 890.77 L776.43 886.29 L766.24 855.73 L768.11 851.21 L807.25 836.89 Z"
      /><path d="M807.25 836.89 L828.26 866.42 L810.8 890.77 L776.43 886.29 L766.24 855.73 L768.11 851.21 L807.25 836.89 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1334.9301 39.94 L1298.71 36.45 L1285.28 51.19 L1293.42 82.99 L1295.78 83.87 L1339.8101 69.47 L1341.35 47.64 L1334.9301 39.94 Z"
      /><path d="M1334.9301 39.94 L1298.71 36.45 L1285.28 51.19 L1293.42 82.99 L1295.78 83.87 L1339.8101 69.47 L1341.35 47.64 L1334.9301 39.94 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M899.26 303.45 L919.47 307.06 L933.34 328.14 L929.17 343.39 L895.63 356.02 L874.05 341.76 L873.73 333.95 L899.26 303.45 Z"
      /><path d="M899.26 303.45 L919.47 307.06 L933.34 328.14 L929.17 343.39 L895.63 356.02 L874.05 341.76 L873.73 333.95 L899.26 303.45 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1551.5 0 L1598 0 L1599.71 40.65 L1584.79 54.22 L1550.34 39 L1551.5 0 Z"
      /><path d="M1551.5 0 L1598 0 L1599.71 40.65 L1584.79 54.22 L1550.34 39 L1551.5 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1299.6 236.39 L1297.21 266.75 L1264.74 269.07 L1242.95 231.69 L1267.59 215.7 L1299.6 236.39 Z"
      /><path d="M1299.6 236.39 L1297.21 266.75 L1264.74 269.07 L1242.95 231.69 L1267.59 215.7 L1299.6 236.39 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M937.75 128.48 L907.38 121.6 L893.5 134.16 L891.65 146.96 L916.46 167.32 L943.1 152.5 L937.75 128.48 Z"
      /><path d="M937.75 128.48 L907.38 121.6 L893.5 134.16 L891.65 146.96 L916.46 167.32 L943.1 152.5 L937.75 128.48 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M958.56 776.81 L937.77 740.62 L910.74 750.48 L907.04 789.93 L941.32 796.47 L958.56 776.81 Z"
      /><path d="M958.56 776.81 L937.77 740.62 L910.74 750.48 L907.04 789.93 L941.32 796.47 L958.56 776.81 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1502.23 223.75 L1481.5 201.87 L1453.1801 209.61 L1448.89 225.56 L1479.9301 255.26 L1492.97 250.46 L1502.23 223.75 Z"
      /><path d="M1502.23 223.75 L1481.5 201.87 L1453.1801 209.61 L1448.89 225.56 L1479.9301 255.26 L1492.97 250.46 L1502.23 223.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1575.04 211.24 L1601.74 212.06 L1615.63 237.32 L1601.08 257.8 L1576.13 252.07 L1567.4399 219.02 L1575.04 211.24 Z"
      /><path d="M1575.04 211.24 L1601.74 212.06 L1615.63 237.32 L1601.08 257.8 L1576.13 252.07 L1567.4399 219.02 L1575.04 211.24 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M388.46 584.77 L347.82 574.24 L330.37 608.73 L340.59 630.61 L363.82 632.41 L389.85 604.2 L388.46 584.77 Z"
      /><path d="M388.46 584.77 L347.82 574.24 L330.37 608.73 L340.59 630.61 L363.82 632.41 L389.85 604.2 L388.46 584.77 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1725.12 219.18 L1697.9 243.59 L1682.29 236.85 L1677.91 193.05 L1707.4 184.11 L1725.12 219.18 Z"
      /><path d="M1725.12 219.18 L1697.9 243.59 L1682.29 236.85 L1677.91 193.05 L1707.4 184.11 L1725.12 219.18 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1715.5699 622.87 L1700.05 648.99 L1679.0699 648.03 L1669.3 622.55 L1694.23 600.99 L1715.5699 622.87 Z"
      /><path d="M1715.5699 622.87 L1700.05 648.99 L1679.0699 648.03 L1669.3 622.55 L1694.23 600.99 L1715.5699 622.87 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1035.88 37.08 L1000.83 28.15 L982.91 54.64 L1013.07 76.53 L1040.23 50.28 L1035.88 37.08 Z"
      /><path d="M1035.88 37.08 L1000.83 28.15 L982.91 54.64 L1013.07 76.53 L1040.23 50.28 L1035.88 37.08 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M225.9 163.84 L207.23 156.78 L178.73 181.27 L180.14 196.88 L209.89 216.96 L218.3 211.75 L226.08 164.11 L225.9 163.84 Z"
      /><path d="M225.9 163.84 L207.23 156.78 L178.73 181.27 L180.14 196.88 L209.89 216.96 L218.3 211.75 L226.08 164.11 L225.9 163.84 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1165.6 0 L1167.66 33.83 L1180.3199 40.3 L1211.52 21.38 L1214.8 0 L1165.6 0 Z"
      /><path d="M1165.6 0 L1167.66 33.83 L1180.3199 40.3 L1211.52 21.38 L1214.8 0 L1165.6 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1124.12 369.29 L1112.77 368.32 L1086.6 406.73 L1111.52 433.34 L1136.02 424.95 L1145 393.03 L1124.12 369.29 Z"
      /><path d="M1124.12 369.29 L1112.77 368.32 L1086.6 406.73 L1111.52 433.34 L1136.02 424.95 L1145 393.03 L1124.12 369.29 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1370.8101 585.77 L1391.3 602.91 L1377.53 629.47 L1338.09 626.6 L1336.17 598.08 L1370.8101 585.77 Z"
      /><path d="M1370.8101 585.77 L1391.3 602.91 L1377.53 629.47 L1338.09 626.6 L1336.17 598.08 L1370.8101 585.77 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M424.42 105.93 L439.04 147.17 L430.66 165.82 L394.2 157.52 L383.97 117.24 L397.34 106.07 L424.42 105.93 Z"
      /><path d="M424.42 105.93 L439.04 147.17 L430.66 165.82 L394.2 157.52 L383.97 117.24 L397.34 106.07 L424.42 105.93 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1061.53 926.05 L1044.84 905.86 L1010.04 907.21 L1003.63 913.93 L1011.13 953.43 L1035.45 961.97 L1061.53 926.05 Z"
      /><path d="M1061.53 926.05 L1044.84 905.86 L1010.04 907.21 L1003.63 913.93 L1011.13 953.43 L1035.45 961.97 L1061.53 926.05 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M197.79 565.9 L179.7 609.15 L222.48 623.62 L231.39 619.33 L237.33 579.2 L197.79 565.9 Z"
      /><path d="M197.79 565.9 L179.7 609.15 L222.48 623.62 L231.39 619.33 L237.33 579.2 L197.79 565.9 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M527.88 959.67 L511.02 987.63 L489.98 985.88 L469.09 955.65 L469.39 952.48 L509.13 932.56 L527.88 959.67 Z"
      /><path d="M527.88 959.67 L511.02 987.63 L489.98 985.88 L469.09 955.65 L469.39 952.48 L509.13 932.56 L527.88 959.67 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1859.1801 1024.62 L1836.99 1019.63 L1811.1801 1036.6 L1811 1080 L1861.1 1080 L1868.71 1046.59 L1859.1801 1024.62 Z"
      /><path d="M1859.1801 1024.62 L1836.99 1019.63 L1811.1801 1036.6 L1811 1080 L1861.1 1080 L1868.71 1046.59 L1859.1801 1024.62 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1217.38 920.1 L1236.63 931.17 L1236.1801 961.05 L1218.05 972.94 L1186.78 954.04 L1187.84 934.68 L1217.38 920.1 Z"
      /><path d="M1217.38 920.1 L1236.63 931.17 L1236.1801 961.05 L1218.05 972.94 L1186.78 954.04 L1187.84 934.68 L1217.38 920.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1416.72 816.25 L1392.92 858.01 L1391.61 858.61 L1361.03 836.66 L1363.77 805.77 L1380.71 792.56 L1389.11 792.48 L1416.72 816.25 Z"
      /><path d="M1416.72 816.25 L1392.92 858.01 L1391.61 858.61 L1361.03 836.66 L1363.77 805.77 L1380.71 792.56 L1389.11 792.48 L1416.72 816.25 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1754.55 764.79 L1716.54 762.15 L1713.1 765.22 L1712.6 808.1 L1732.9301 817.04 L1759.08 800.59 L1754.55 764.79 Z"
      /><path d="M1754.55 764.79 L1716.54 762.15 L1713.1 765.22 L1712.6 808.1 L1732.9301 817.04 L1759.08 800.59 L1754.55 764.79 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M279.8 154.9 L317.62 169.04 L316.01 187.35 L288.99 201.16 L265.5 187.6 L262.87 177.8 L279.8 154.9 Z"
      /><path d="M279.8 154.9 L317.62 169.04 L316.01 187.35 L288.99 201.16 L265.5 187.6 L262.87 177.8 L279.8 154.9 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M776.43 886.29 L810.8 890.77 L820.83 918.6 L812.13 935.41 L773 939.25 L761.68 907.08 L776.43 886.29 Z"
      /><path d="M776.43 886.29 L810.8 890.77 L820.83 918.6 L812.13 935.41 L773 939.25 L761.68 907.08 L776.43 886.29 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1153.99 334.45 L1136.0699 308.24 L1101.7 317.62 L1094.63 349.46 L1112.77 368.32 L1124.12 369.29 L1153.99 334.45 Z"
      /><path d="M1153.99 334.45 L1136.0699 308.24 L1101.7 317.62 L1094.63 349.46 L1112.77 368.32 L1124.12 369.29 L1153.99 334.45 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1528.27 713.07 L1527.38 747.7 L1490.74 756.74 L1476.84 732.65 L1483.0601 713.66 L1497.4399 704.62 L1528.27 713.07 Z"
      /><path d="M1528.27 713.07 L1527.38 747.7 L1490.74 756.74 L1476.84 732.65 L1483.0601 713.66 L1497.4399 704.62 L1528.27 713.07 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1103.6899 456.55 L1117 478.95 L1099.58 511.37 L1082.67 513.1 L1059.5 489.59 L1063.16 463.82 L1103.6899 456.55 Z"
      /><path d="M1103.6899 456.55 L1117 478.95 L1099.58 511.37 L1082.67 513.1 L1059.5 489.59 L1063.16 463.82 L1103.6899 456.55 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M56.62 654.41 L51.3 659.49 L0 659.2 L0 607.1 L43.46 603.18 L56.62 654.41 Z"
      /><path d="M56.62 654.41 L51.3 659.49 L0 659.2 L0 607.1 L43.46 603.18 L56.62 654.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1102.67 667.12 L1069.74 649.45 L1050.76 657.78 L1047.13 701.58 L1049.04 704.4 L1090.24 701.39 L1104.9399 675.44 L1102.67 667.12 Z"
      /><path d="M1102.67 667.12 L1069.74 649.45 L1050.76 657.78 L1047.13 701.58 L1049.04 704.4 L1090.24 701.39 L1104.9399 675.44 L1102.67 667.12 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M1920 415.8 L1874.17 403.56 L1869.71 405.13 L1862.89 430.23 L1877.5601 452.64 L1920 443.7 L1920 415.8 Z"
      /><path d="M1920 415.8 L1874.17 403.56 L1869.71 405.13 L1862.89 430.23 L1877.5601 452.64 L1920 443.7 L1920 415.8 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1285.28 51.19 L1255.8 43.42 L1235.37 55.6 L1234.0601 58.59 L1235.92 76 L1254.01 95.75 L1270.09 97.69 L1293.42 82.99 L1285.28 51.19 Z"
      /><path d="M1285.28 51.19 L1255.8 43.42 L1235.37 55.6 L1234.0601 58.59 L1235.92 76 L1254.01 95.75 L1270.09 97.69 L1293.42 82.99 L1285.28 51.19 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1005 1080 L982.75 1030.75 L968.54 1031.25 L948.85 1052.3199 L952 1080 L1005 1080 Z"
      /><path d="M1005 1080 L982.75 1030.75 L968.54 1031.25 L948.85 1052.3199 L952 1080 L1005 1080 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1230.13 831.05 L1227.92 828.96 L1189.52 834.64 L1183.55 849 L1196.05 880.8 L1213.75 886.6 L1233.39 874.91 L1230.13 831.05 Z"
      /><path d="M1230.13 831.05 L1227.92 828.96 L1189.52 834.64 L1183.55 849 L1196.05 880.8 L1213.75 886.6 L1233.39 874.91 L1230.13 831.05 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1237.0699 690.06 L1259.28 711.73 L1254.46 734.96 L1221.15 747.73 L1196.42 721.82 L1204.77 697.74 L1237.0699 690.06 Z"
      /><path d="M1237.0699 690.06 L1259.28 711.73 L1254.46 734.96 L1221.15 747.73 L1196.42 721.82 L1204.77 697.74 L1237.0699 690.06 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M941.18 993.83 L940.97 996.41 L917.04 1020.82 L887.54 1012.41 L878.6 993.78 L915.26 970.5 L941.18 993.83 Z"
      /><path d="M941.18 993.83 L940.97 996.41 L917.04 1020.82 L887.54 1012.41 L878.6 993.78 L915.26 970.5 L941.18 993.83 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M654.94 298.62 L621.86 262.32 L615.46 263.35 L590.12 305.37 L612.88 329.98 L617.62 331.02 L652.81 310.23 L654.94 298.62 Z"
      /><path d="M654.94 298.62 L621.86 262.32 L615.46 263.35 L590.12 305.37 L612.88 329.98 L617.62 331.02 L652.81 310.23 L654.94 298.62 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M262.07 313.98 L234.78 304.04 L213.77 315.16 L208.74 341.01 L233.15 359.58 L251.75 355.45 L263.24 316.12 L262.07 313.98 Z"
      /><path d="M262.07 313.98 L234.78 304.04 L213.77 315.16 L208.74 341.01 L233.15 359.58 L251.75 355.45 L263.24 316.12 L262.07 313.98 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1418.89 564.96 L1403.91 540.07 L1369.59 557.15 L1370.8101 585.77 L1391.3 602.91 L1398.9399 601.52 L1418.89 564.96 Z"
      /><path d="M1418.89 564.96 L1403.91 540.07 L1369.59 557.15 L1370.8101 585.77 L1391.3 602.91 L1398.9399 601.52 L1418.89 564.96 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M836.94 529.63 L869.15 542.3 L873.76 551.83 L848.15 588.48 L842.95 589.17 L813.79 557.64 L815.8 545.16 L836.94 529.63 Z"
      /><path d="M836.94 529.63 L869.15 542.3 L873.76 551.83 L848.15 588.48 L842.95 589.17 L813.79 557.64 L815.8 545.16 L836.94 529.63 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M730.61 1039.0601 L703.79 1028.97 L692.2 1035.17 L690.9 1080 L732.6 1080 L730.61 1039.0601 Z"
      /><path d="M730.61 1039.0601 L703.79 1028.97 L692.2 1035.17 L690.9 1080 L732.6 1080 L730.61 1039.0601 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1055.74 873.61 L1044.84 905.86 L1010.04 907.21 L1004.14 863.84 L1033.1801 852.13 L1055.74 873.61 Z"
      /><path d="M1055.74 873.61 L1044.84 905.86 L1010.04 907.21 L1004.14 863.84 L1033.1801 852.13 L1055.74 873.61 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1254.01 95.75 L1232.78 128.19 L1216.8 129.24 L1203.64 100.69 L1235.92 76 L1254.01 95.75 Z"
      /><path d="M1254.01 95.75 L1232.78 128.19 L1216.8 129.24 L1203.64 100.69 L1235.92 76 L1254.01 95.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M561.03 171.49 L583.65 206.15 L575.69 224.19 L522.29 218.74 L523.42 187.06 L561.03 171.49 Z"
      /><path d="M561.03 171.49 L583.65 206.15 L575.69 224.19 L522.29 218.74 L523.42 187.06 L561.03 171.49 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M790.8 115.41 L766.67 103.77 L746.52 113.84 L760.31 156.27 L771.29 159.63 L795.5 129.14 L790.8 115.41 Z"
      /><path d="M790.8 115.41 L766.67 103.77 L746.52 113.84 L760.31 156.27 L771.29 159.63 L795.5 129.14 L790.8 115.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1601.1801 722.35 L1579.21 727.43 L1570.73 751.87 L1584.99 770.94 L1614.12 771.64 L1623.71 761.78 L1624.79 742.97 L1601.1801 722.35 Z"
      /><path d="M1601.1801 722.35 L1579.21 727.43 L1570.73 751.87 L1584.99 770.94 L1614.12 771.64 L1623.71 761.78 L1624.79 742.97 L1601.1801 722.35 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M102.48 88.92 L102.67 88.94 L125.95 116.48 L122.77 131.98 L100.82 143.49 L76.99 112.21 L102.48 88.92 Z"
      /><path d="M102.48 88.92 L102.67 88.94 L125.95 116.48 L122.77 131.98 L100.82 143.49 L76.99 112.21 L102.48 88.92 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1035.45 961.97 L1011.13 953.43 L981.79 972.02 L1001.66 1012.65 L1020.45 1013.34 L1042.24 976.05 L1035.45 961.97 Z"
      /><path d="M1035.45 961.97 L1011.13 953.43 L981.79 972.02 L1001.66 1012.65 L1020.45 1013.34 L1042.24 976.05 L1035.45 961.97 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1068 601.08 L1077.3199 612.16 L1069.74 649.45 L1050.76 657.78 L1028.23 645.64 L1022.44 621.49 L1040.74 599.75 L1068 601.08 Z"
      /><path d="M1068 601.08 L1077.3199 612.16 L1069.74 649.45 L1050.76 657.78 L1028.23 645.64 L1022.44 621.49 L1040.74 599.75 L1068 601.08 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M657.94 1003.58 L665.55 1028.35 L649.26 1044.41 L613.74 1037.5699 L610.14 1032.3101 L623.12 996.34 L657.94 1003.58 Z"
      /><path d="M657.94 1003.58 L665.55 1028.35 L649.26 1044.41 L613.74 1037.5699 L610.14 1032.3101 L623.12 996.34 L657.94 1003.58 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M468.84 449.46 L448.8 475.17 L466.73 500.79 L487.61 501.21 L500.61 477.86 L485.93 451.89 L468.84 449.46 Z"
      /><path d="M468.84 449.46 L448.8 475.17 L466.73 500.79 L487.61 501.21 L500.61 477.86 L485.93 451.89 L468.84 449.46 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M396.56 1027.0601 L429.65 1042 L432.6 1080 L377.8 1080 L376.77 1045.8199 L396.56 1027.0601 Z"
      /><path d="M396.56 1027.0601 L429.65 1042 L432.6 1080 L377.8 1080 L376.77 1045.8199 L396.56 1027.0601 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1567.4399 219.02 L1537.74 219.4 L1535.54 269.29 L1550.95 272.79 L1576.13 252.07 L1567.4399 219.02 Z"
      /><path d="M1567.4399 219.02 L1537.74 219.4 L1535.54 269.29 L1550.95 272.79 L1576.13 252.07 L1567.4399 219.02 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M359.56 738.1 L342.34 701.86 L307.44 711.48 L308.05 751.12 L316.62 760.06 L346.66 757.94 L359.56 738.1 Z"
      /><path d="M359.56 738.1 L342.34 701.86 L307.44 711.48 L308.05 751.12 L316.62 760.06 L346.66 757.94 L359.56 738.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M621.16 470.64 L639.61 476.76 L650.16 522.05 L647.28 526.42 L608.37 528.57 L603.74 479.96 L621.16 470.64 Z"
      /><path d="M621.16 470.64 L639.61 476.76 L650.16 522.05 L647.28 526.42 L608.37 528.57 L603.74 479.96 L621.16 470.64 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1641.65 517.77 L1619.76 546.25 L1602.1801 542.44 L1587.55 521.9 L1598.05 491.93 L1623.87 482.73 L1641.65 517.77 Z"
      /><path d="M1641.65 517.77 L1619.76 546.25 L1602.1801 542.44 L1587.55 521.9 L1598.05 491.93 L1623.87 482.73 L1641.65 517.77 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M426.41 474.82 L448.8 475.17 L466.73 500.79 L441.53 533.45 L435.72 531.43 L415.2 498.51 L426.41 474.82 Z"
      /><path d="M426.41 474.82 L448.8 475.17 L466.73 500.79 L441.53 533.45 L435.72 531.43 L415.2 498.51 L426.41 474.82 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1833.6801 681.29 L1812.64 651.51 L1793.23 652.88 L1777.33 678.61 L1792.45 707.66 L1809.04 711.71 L1826.96 701.99 L1833.6801 681.29 Z"
      /><path d="M1833.6801 681.29 L1812.64 651.51 L1793.23 652.88 L1777.33 678.61 L1792.45 707.66 L1809.04 711.71 L1826.96 701.99 L1833.6801 681.29 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M210.58 951.25 L244.09 968.82 L246.3 991.33 L219.29 1017.45 L182.37 991.96 L188.17 965.95 L210.58 951.25 Z"
      /><path d="M210.58 951.25 L244.09 968.82 L246.3 991.33 L219.29 1017.45 L182.37 991.96 L188.17 965.95 L210.58 951.25 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1814.38 231.44 L1797.89 227.47 L1773.99 253.27 L1786.64 275.57 L1821.96 276.34 L1829.28 262.87 L1814.38 231.44 Z"
      /><path d="M1814.38 231.44 L1797.89 227.47 L1773.99 253.27 L1786.64 275.57 L1821.96 276.34 L1829.28 262.87 L1814.38 231.44 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M198.32 86.07 L184.03 81.23 L159.05 96.42 L158.14 99.31 L171.68 131.44 L196.81 135.13 L209.93 112.07 L198.32 86.07 Z"
      /><path d="M198.32 86.07 L184.03 81.23 L159.05 96.42 L158.14 99.31 L171.68 131.44 L196.81 135.13 L209.93 112.07 L198.32 86.07 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1332.53 633.94 L1336.8101 668.87 L1293.39 675.43 L1281.67 656.51 L1293.45 631.48 L1332.53 633.94 Z"
      /><path d="M1332.53 633.94 L1336.8101 668.87 L1293.39 675.43 L1281.67 656.51 L1293.45 631.48 L1332.53 633.94 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1347.55 928.47 L1332.73 936.85 L1328.4 974.22 L1365.36 991.44 L1372.8199 987.48 L1387.1 951.67 L1382.79 941.89 L1347.55 928.47 Z"
      /><path d="M1347.55 928.47 L1332.73 936.85 L1328.4 974.22 L1365.36 991.44 L1372.8199 987.48 L1387.1 951.67 L1382.79 941.89 L1347.55 928.47 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1920 242.7 L1873.87 264.45 L1876.25 296.22 L1889.04 306.35 L1920 304.9 L1920 242.7 Z"
      /><path d="M1920 242.7 L1873.87 264.45 L1876.25 296.22 L1889.04 306.35 L1920 304.9 L1920 242.7 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1715.4399 722.56 L1699.78 713.58 L1669.97 735.46 L1676 762.72 L1713.1 765.22 L1716.54 762.15 L1715.4399 722.56 Z"
      /><path d="M1715.4399 722.56 L1699.78 713.58 L1669.97 735.46 L1676 762.72 L1713.1 765.22 L1716.54 762.15 L1715.4399 722.56 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M571.96 599.49 L540.07 613.4 L549.13 651.42 L584.23 646.89 L593.45 627.44 L571.96 599.49 Z"
      /><path d="M571.96 599.49 L540.07 613.4 L549.13 651.42 L584.23 646.89 L593.45 627.44 L571.96 599.49 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1858.49 144.85 L1804.3199 118.91 L1797.21 125.32 L1791.29 146.19 L1812.2 175.39 L1825.73 176.97 L1858.49 144.87 L1858.49 144.85 Z"
      /><path d="M1858.49 144.85 L1804.3199 118.91 L1797.21 125.32 L1791.29 146.19 L1812.2 175.39 L1825.73 176.97 L1858.49 144.87 L1858.49 144.85 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1631.48 99.71 L1612.4301 132.81 L1620.46 151.82 L1657.4399 153.61 L1674.46 131.47 L1672.52 121.11 L1631.48 99.71 Z"
      /><path d="M1631.48 99.71 L1612.4301 132.81 L1620.46 151.82 L1657.4399 153.61 L1674.46 131.47 L1672.52 121.11 L1631.48 99.71 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M812.4 36.93 L781.96 35.92 L764.15 58.04 L772.12 71.31 L815.99 75.57 L815.66 40.29 L812.4 36.93 Z"
      /><path d="M812.4 36.93 L781.96 35.92 L764.15 58.04 L772.12 71.31 L815.99 75.57 L815.66 40.29 L812.4 36.93 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M455.54 767.65 L454.1 795.44 L416.42 807.34 L398.64 783.9 L407.52 758.11 L439.41 752.39 L455.54 767.65 Z"
      /><path d="M455.54 767.65 L454.1 795.44 L416.42 807.34 L398.64 783.9 L407.52 758.11 L439.41 752.39 L455.54 767.65 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M108.6 517.2 L129.38 523.35 L142.31 558.6 L135.95 570.82 L95.5 576.8 L81.57 536.16 L108.6 517.2 Z"
      /><path d="M108.6 517.2 L129.38 523.35 L142.31 558.6 L135.95 570.82 L95.5 576.8 L81.57 536.16 L108.6 517.2 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1620.66 807.62 L1600.45 820.23 L1601.5 854.96 L1634.14 861.21 L1648.99 842.56 L1639.54 813.74 L1620.66 807.62 Z"
      /><path d="M1620.66 807.62 L1600.45 820.23 L1601.5 854.96 L1634.14 861.21 L1648.99 842.56 L1639.54 813.74 L1620.66 807.62 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M560.13 805.41 L564.3 812.76 L560.34 838.95 L523.02 855.61 L514.29 851.73 L515.12 813.83 L560.13 805.41 Z"
      /><path d="M560.13 805.41 L564.3 812.76 L560.34 838.95 L523.02 855.61 L514.29 851.73 L515.12 813.83 L560.13 805.41 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M179.7 609.15 L222.48 623.62 L209.42 666.77 L205.02 668.1 L173.21 653.57 L177.28 610.31 L179.7 609.15 Z"
      /><path d="M179.7 609.15 L222.48 623.62 L209.42 666.77 L205.02 668.1 L173.21 653.57 L177.28 610.31 L179.7 609.15 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M650.7 0 L648.81 42.16 L642.61 46.45 L599.97 40.53 L596.6 0 L650.7 0 Z"
      /><path d="M650.7 0 L648.81 42.16 L642.61 46.45 L599.97 40.53 L596.6 0 L650.7 0 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1534.38 663.82 L1571.74 667.54 L1577.45 674.82 L1562.88 708.94 L1534.63 708.33 L1534.38 663.82 Z"
      /><path d="M1534.38 663.82 L1571.74 667.54 L1577.45 674.82 L1562.88 708.94 L1534.63 708.33 L1534.38 663.82 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1641.1899 955.33 L1655.11 957.31 L1677.77 986.89 L1668.58 1021.83 L1625.95 1023.34 L1612.27 1003.45 L1619.58 968.91 L1641.1899 955.33 Z"
      /><path d="M1641.1899 955.33 L1655.11 957.31 L1677.77 986.89 L1668.58 1021.83 L1625.95 1023.34 L1612.27 1003.45 L1619.58 968.91 L1641.1899 955.33 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1517.55 836.36 L1485.6801 850.72 L1486.61 875.81 L1503.55 889.62 L1530.03 879.33 L1530.29 843.66 L1517.55 836.36 Z"
      /><path d="M1517.55 836.36 L1485.6801 850.72 L1486.61 875.81 L1503.55 889.62 L1530.03 879.33 L1530.29 843.66 L1517.55 836.36 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1325.74 474.37 L1323.37 473.87 L1292.21 490.02 L1289.8199 515.82 L1304.74 528.4 L1343.39 515.17 L1325.74 474.37 Z"
      /><path d="M1325.74 474.37 L1323.37 473.87 L1292.21 490.02 L1289.8199 515.82 L1304.74 528.4 L1343.39 515.17 L1325.74 474.37 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1040.23 50.28 L1063.12 62.24 L1063.17 84.42 L1041.99 101.03 L1014.8 87.25 L1013.07 76.53 L1040.23 50.28 Z"
      /><path d="M1040.23 50.28 L1063.12 62.24 L1063.17 84.42 L1041.99 101.03 L1014.8 87.25 L1013.07 76.53 L1040.23 50.28 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M642.61 46.45 L599.97 40.53 L592.17 49.19 L603.85 93.07 L634.78 93.96 L642.61 46.45 Z"
      /><path d="M642.61 46.45 L599.97 40.53 L592.17 49.19 L603.85 93.07 L634.78 93.96 L642.61 46.45 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M922.97 38.36 L919.69 53.37 L891.85 60.73 L874.04 43.79 L898.41 12.65 L922.97 38.36 Z"
      /><path d="M922.97 38.36 L919.69 53.37 L891.85 60.73 L874.04 43.79 L898.41 12.65 L922.97 38.36 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M772.72 1036.89 L753.92 1025.98 L730.61 1039.0601 L732.6 1080 L769.3 1080 L772.72 1036.89 Z"
      /><path d="M772.72 1036.89 L753.92 1025.98 L730.61 1039.0601 L732.6 1080 L769.3 1080 L772.72 1036.89 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1092.49 851.62 L1084.63 868.16 L1055.74 873.61 L1033.1801 852.13 L1038.8 827.94 L1076.67 818.33 L1092.49 851.62 Z"
      /><path d="M1092.49 851.62 L1084.63 868.16 L1055.74 873.61 L1033.1801 852.13 L1038.8 827.94 L1076.67 818.33 L1092.49 851.62 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M1763.97 730.85 L1739.62 713.88 L1715.4399 722.56 L1716.54 762.15 L1754.55 764.79 L1765.52 753.44 L1763.97 730.85 Z"
      /><path d="M1763.97 730.85 L1739.62 713.88 L1715.4399 722.56 L1716.54 762.15 L1754.55 764.79 L1765.52 753.44 L1763.97 730.85 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1566 807.77 L1552.8 836.35 L1530.29 843.66 L1517.55 836.36 L1510.1 802.19 L1535.9301 789.34 L1566 807.77 Z"
      /><path d="M1566 807.77 L1552.8 836.35 L1530.29 843.66 L1517.55 836.36 L1510.1 802.19 L1535.9301 789.34 L1566 807.77 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M282.39 453.74 L328.89 469.16 L322.11 502.54 L312.66 508.28 L274.19 494.38 L268.31 469.82 L282.39 453.74 Z"
      /><path d="M282.39 453.74 L328.89 469.16 L322.11 502.54 L312.66 508.28 L274.19 494.38 L268.31 469.82 L282.39 453.74 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1765.0601 197.15 L1786.53 202.69 L1797.89 227.47 L1773.99 253.27 L1755.76 250.33 L1742.04 222.3 L1765.0601 197.15 Z"
      /><path d="M1765.0601 197.15 L1786.53 202.69 L1797.89 227.47 L1773.99 253.27 L1755.76 250.33 L1742.04 222.3 L1765.0601 197.15 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M776.43 886.29 L766.24 855.73 L714.68 866.34 L728.43 904.21 L761.68 907.08 L776.43 886.29 Z"
      /><path d="M776.43 886.29 L766.24 855.73 L714.68 866.34 L728.43 904.21 L761.68 907.08 L776.43 886.29 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1624.0601 329.35 L1619 339.09 L1585.96 348.11 L1563.17 322.56 L1569.7 302.94 L1607.84 291.38 L1624.0601 329.35 Z"
      /><path d="M1624.0601 329.35 L1619 339.09 L1585.96 348.11 L1563.17 322.56 L1569.7 302.94 L1607.84 291.38 L1624.0601 329.35 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M151.11 162.7 L178.73 181.27 L180.14 196.88 L154.2 216.22 L139 210.26 L130.63 181.81 L151.11 162.7 Z"
      /><path d="M151.11 162.7 L178.73 181.27 L180.14 196.88 L154.2 216.22 L139 210.26 L130.63 181.81 L151.11 162.7 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M612.88 329.98 L575.42 369.03 L575.53 370.92 L601.49 390.81 L636.76 371.08 L617.62 331.02 L612.88 329.98 Z"
      /><path d="M612.88 329.98 L575.42 369.03 L575.53 370.92 L601.49 390.81 L636.76 371.08 L617.62 331.02 L612.88 329.98 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M414.21 913.51 L425.63 928.74 L409.87 960.75 L379.2 954.88 L372.15 919.63 L414.21 913.51 Z"
      /><path d="M414.21 913.51 L425.63 928.74 L409.87 960.75 L379.2 954.88 L372.15 919.63 L414.21 913.51 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1766.85 357.8 L1748.77 351.56 L1722.5699 367.48 L1719.8101 387.22 L1750.48 411.22 L1774.8101 388.99 L1766.85 357.8 Z"
      /><path d="M1766.85 357.8 L1748.77 351.56 L1722.5699 367.48 L1719.8101 387.22 L1750.48 411.22 L1774.8101 388.99 L1766.85 357.8 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M164.2 303.86 L139.51 285.26 L114.08 297.04 L111.6 323.27 L132.36 340.13 L160.07 327.09 L164.2 303.86 Z"
      /><path d="M164.2 303.86 L139.51 285.26 L114.08 297.04 L111.6 323.27 L132.36 340.13 L160.07 327.09 L164.2 303.86 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M764.15 58.04 L738.99 52.64 L733.4 55.09 L721.06 94.31 L735.51 111.62 L746.52 113.84 L766.67 103.77 L772.12 71.31 L764.15 58.04 Z"
      /><path d="M764.15 58.04 L738.99 52.64 L733.4 55.09 L721.06 94.31 L735.51 111.62 L746.52 113.84 L766.67 103.77 L772.12 71.31 L764.15 58.04 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M330.37 608.73 L340.59 630.61 L325.12 653.07 L305.94 656.28 L277.53 626.61 L290.51 600.39 L330.37 608.73 Z"
      /><path d="M330.37 608.73 L340.59 630.61 L325.12 653.07 L305.94 656.28 L277.53 626.61 L290.51 600.39 L330.37 608.73 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1871.85 846.1 L1907.65 874.15 L1871.54 905.64 L1849.7 883.07 L1855.99 849.83 L1871.85 846.1 Z"
      /><path d="M1871.85 846.1 L1907.65 874.15 L1871.54 905.64 L1849.7 883.07 L1855.99 849.83 L1871.85 846.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M218.3 211.75 L209.89 216.96 L209.08 220.61 L227.75 263.29 L231.31 264.78 L251.51 257.39 L259.4 235.26 L245.91 214.63 L218.3 211.75 Z"
      /><path d="M218.3 211.75 L209.89 216.96 L209.08 220.61 L227.75 263.29 L231.31 264.78 L251.51 257.39 L259.4 235.26 L245.91 214.63 L218.3 211.75 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M719.69 431.88 L712.24 461.71 L681.1 471.06 L668.51 463.4 L666.46 433.01 L700.52 417.35 L719.69 431.88 Z"
      /><path d="M719.69 431.88 L712.24 461.71 L681.1 471.06 L668.51 463.4 L666.46 433.01 L700.52 417.35 L719.69 431.88 Z" style="fill:rgb(23,201,0); stroke:none;"
      /><path style="fill:none;" d="M1709.85 928.62 L1725.75 972.5 L1724.85 974.55 L1677.77 986.89 L1655.11 957.31 L1686.6801 923.82 L1709.85 928.62 Z"
      /><path d="M1709.85 928.62 L1725.75 972.5 L1724.85 974.55 L1677.77 986.89 L1655.11 957.31 L1686.6801 923.82 L1709.85 928.62 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1640.3199 658.58 L1668.29 660.2 L1674.28 687.65 L1647.64 702.72 L1634.17 693.12 L1640.3199 658.58 Z"
      /><path d="M1640.3199 658.58 L1668.29 660.2 L1674.28 687.65 L1647.64 702.72 L1634.17 693.12 L1640.3199 658.58 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1353.52 268.67 L1378.1801 270.19 L1397.41 293.45 L1386.1801 326.64 L1370.6801 333.49 L1342.34 320.92 L1350.8 270.86 L1353.52 268.67 Z"
      /><path d="M1353.52 268.67 L1378.1801 270.19 L1397.41 293.45 L1386.1801 326.64 L1370.6801 333.49 L1342.34 320.92 L1350.8 270.86 L1353.52 268.67 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M205.02 668.1 L185.83 710.79 L163.42 709.4 L146.23 666.74 L173.21 653.57 L205.02 668.1 Z"
      /><path d="M205.02 668.1 L185.83 710.79 L163.42 709.4 L146.23 666.74 L173.21 653.57 L205.02 668.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1314.8 360.56 L1321.41 375.04 L1301.5 413.86 L1256.78 379.3 L1276.92 352.59 L1314.8 360.56 Z"
      /><path d="M1314.8 360.56 L1321.41 375.04 L1301.5 413.86 L1256.78 379.3 L1276.92 352.59 L1314.8 360.56 Z" style="fill:rgb(35,189,0); stroke:none;"
      /><path style="fill:none;" d="M134.03 52.18 L132.33 67.23 L102.67 88.94 L102.48 88.92 L81.71 62.36 L84.8 46.12 L114.54 37.01 L134.03 52.18 Z"
      /><path d="M134.03 52.18 L132.33 67.23 L102.67 88.94 L102.48 88.92 L81.71 62.36 L84.8 46.12 L114.54 37.01 L134.03 52.18 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1844.87 345.48 L1815.33 354.62 L1811.33 396.03 L1853 391.78 L1853 350.38 L1844.87 345.48 Z"
      /><path d="M1844.87 345.48 L1815.33 354.62 L1811.33 396.03 L1853 391.78 L1853 350.38 L1844.87 345.48 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1020.75 343.39 L1008.16 332.35 L982.07 334.86 L968.88 372.04 L975.92 380.31 L1013.3 380.96 L1020.75 343.39 Z"
      /><path d="M1020.75 343.39 L1008.16 332.35 L982.07 334.86 L968.88 372.04 L975.92 380.31 L1013.3 380.96 L1020.75 343.39 Z" style="fill:rgb(11,213,0); stroke:none;"
      /><path style="fill:none;" d="M551.47 959.1 L568.12 993.83 L565.97 999.27 L524.32 1007.81 L511.02 987.63 L527.88 959.67 L551.47 959.1 Z"
      /><path d="M551.47 959.1 L568.12 993.83 L565.97 999.27 L524.32 1007.81 L511.02 987.63 L527.88 959.67 L551.47 959.1 Z" style="fill:rgb(0,0,139); stroke:none;"
      /><path style="fill:none;" d="M1407.6899 435.48 L1365.66 422.98 L1359.45 428.61 L1353.6801 457.3 L1386.13 484.95 L1409.78 472.26 L1407.6899 435.48 Z"
      /><path d="M1407.6899 435.48 L1365.66 422.98 L1359.45 428.61 L1353.6801 457.3 L1386.13 484.95 L1409.78 472.26 L1407.6899 435.48 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1407.6899 435.48 L1365.66 422.98 L1359.45 428.61 L1353.6801 457.3 L1386.13 484.95 L1409.78 472.26 L1407.6899 435.48 Z"
      /><path d="M1407.6899 435.48 L1365.66 422.98 L1359.45 428.61 L1353.6801 457.3 L1386.13 484.95 L1409.78 472.26 L1407.6899 435.48 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M955.65 935.97 L921.95 936.04 L914.2 944.68 L915.26 970.5 L941.18 993.83 L973.36 970.28 L955.65 935.97 Z"
      /><path d="M955.65 935.97 L921.95 936.04 L914.2 944.68 L915.26 970.5 L941.18 993.83 L973.36 970.28 L955.65 935.97 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M955.65 935.97 L921.95 936.04 L914.2 944.68 L915.26 970.5 L941.18 993.83 L973.36 970.28 L955.65 935.97 Z"
      /><path d="M955.65 935.97 L921.95 936.04 L914.2 944.68 L915.26 970.5 L941.18 993.83 L973.36 970.28 L955.65 935.97 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M553.34 428.25 L571.04 434.9 L581.12 475.22 L558.18 491.95 L545.94 491.11 L530.85 475.57 L536.26 437.55 L553.34 428.25 Z"
      /><path d="M553.34 428.25 L571.04 434.9 L581.12 475.22 L558.18 491.95 L545.94 491.11 L530.85 475.57 L536.26 437.55 L553.34 428.25 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M553.34 428.25 L571.04 434.9 L581.12 475.22 L558.18 491.95 L545.94 491.11 L530.85 475.57 L536.26 437.55 L553.34 428.25 Z"
      /><path d="M553.34 428.25 L571.04 434.9 L581.12 475.22 L558.18 491.95 L545.94 491.11 L530.85 475.57 L536.26 437.55 L553.34 428.25 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1014.8 87.25 L1041.99 101.03 L1044.47 128.92 L1038 136.43 L990.54 119.73 L989.56 116.82 L1014.8 87.25 Z"
      /><path d="M1014.8 87.25 L1041.99 101.03 L1044.47 128.92 L1038 136.43 L990.54 119.73 L989.56 116.82 L1014.8 87.25 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1142.4 877.99 L1170.33 899.13 L1169.4 917.75 L1133.7 932.8 L1119.51 898.27 L1142.4 877.99 Z"
      /><path d="M1142.4 877.99 L1170.33 899.13 L1169.4 917.75 L1133.7 932.8 L1119.51 898.27 L1142.4 877.99 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1142.4 877.99 L1170.33 899.13 L1169.4 917.75 L1133.7 932.8 L1119.51 898.27 L1142.4 877.99 Z"
      /><path d="M1142.4 877.99 L1170.33 899.13 L1169.4 917.75 L1133.7 932.8 L1119.51 898.27 L1142.4 877.99 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1321.41 375.04 L1301.5 413.86 L1301.76 415.95 L1359.45 428.61 L1365.66 422.98 L1368.3 384.07 L1367.0601 382.52 L1321.41 375.04 Z"
      /><path d="M1321.41 375.04 L1301.5 413.86 L1301.76 415.95 L1359.45 428.61 L1365.66 422.98 L1368.3 384.07 L1367.0601 382.52 L1321.41 375.04 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1321.41 375.04 L1301.5 413.86 L1301.76 415.95 L1359.45 428.61 L1365.66 422.98 L1368.3 384.07 L1367.0601 382.52 L1321.41 375.04 Z"
      /><path d="M1321.41 375.04 L1301.5 413.86 L1301.76 415.95 L1359.45 428.61 L1365.66 422.98 L1368.3 384.07 L1367.0601 382.52 L1321.41 375.04 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1321.41 375.04 L1301.5 413.86 L1301.76 415.95 L1359.45 428.61 L1365.66 422.98 L1368.3 384.07 L1367.0601 382.52 L1321.41 375.04 Z"
      /><path d="M1321.41 375.04 L1301.5 413.86 L1301.76 415.95 L1359.45 428.61 L1365.66 422.98 L1368.3 384.07 L1367.0601 382.52 L1321.41 375.04 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1433.5699 482.78 L1438.78 514.74 L1404.45 537.68 L1380.76 501.69 L1386.13 484.95 L1409.78 472.26 L1433.5699 482.78 Z"
      /><path d="M1433.5699 482.78 L1438.78 514.74 L1404.45 537.68 L1380.76 501.69 L1386.13 484.95 L1409.78 472.26 L1433.5699 482.78 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M549.36 553.89 L546.29 553.73 L523.98 572.82 L527.97 608.02 L540.07 613.4 L571.96 599.49 L575.72 585.44 L549.36 553.89 Z"
      /><path d="M549.36 553.89 L546.29 553.73 L523.98 572.82 L527.97 608.02 L540.07 613.4 L571.96 599.49 L575.72 585.44 L549.36 553.89 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M549.36 553.89 L546.29 553.73 L523.98 572.82 L527.97 608.02 L540.07 613.4 L571.96 599.49 L575.72 585.44 L549.36 553.89 Z"
      /><path d="M549.36 553.89 L546.29 553.73 L523.98 572.82 L527.97 608.02 L540.07 613.4 L571.96 599.49 L575.72 585.44 L549.36 553.89 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M714.68 866.34 L728.43 904.21 L710.43 928.48 L691.35 928.26 L671.4 904.58 L674.67 881.7 L713.54 865.6 L714.68 866.34 Z"
      /><path d="M714.68 866.34 L728.43 904.21 L710.43 928.48 L691.35 928.26 L671.4 904.58 L674.67 881.7 L713.54 865.6 L714.68 866.34 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M671.18 799.59 L640.56 769.98 L617.67 783.67 L616.16 816.42 L660.31 827.04 L666.53 822.38 L671.18 799.59 Z"
      /><path d="M671.18 799.59 L640.56 769.98 L617.67 783.67 L616.16 816.42 L660.31 827.04 L666.53 822.38 L671.18 799.59 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M671.18 799.59 L640.56 769.98 L617.67 783.67 L616.16 816.42 L660.31 827.04 L666.53 822.38 L671.18 799.59 Z"
      /><path d="M671.18 799.59 L640.56 769.98 L617.67 783.67 L616.16 816.42 L660.31 827.04 L666.53 822.38 L671.18 799.59 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M872.35 939.1 L863.13 916.03 L820.83 918.6 L812.13 935.41 L824.35 961.39 L860.07 961.8 L872.35 939.1 Z"
      /><path d="M872.35 939.1 L863.13 916.03 L820.83 918.6 L812.13 935.41 L824.35 961.39 L860.07 961.8 L872.35 939.1 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M872.35 939.1 L863.13 916.03 L820.83 918.6 L812.13 935.41 L824.35 961.39 L860.07 961.8 L872.35 939.1 Z"
      /><path d="M872.35 939.1 L863.13 916.03 L820.83 918.6 L812.13 935.41 L824.35 961.39 L860.07 961.8 L872.35 939.1 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M575.53 370.92 L601.49 390.81 L603.61 419.04 L571.04 434.9 L553.34 428.25 L549.6 393.46 L575.53 370.92 Z"
      /><path d="M575.53 370.92 L601.49 390.81 L603.61 419.04 L571.04 434.9 L553.34 428.25 L549.6 393.46 L575.53 370.92 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M575.53 370.92 L601.49 390.81 L603.61 419.04 L571.04 434.9 L553.34 428.25 L549.6 393.46 L575.53 370.92 Z"
      /><path d="M575.53 370.92 L601.49 390.81 L603.61 419.04 L571.04 434.9 L553.34 428.25 L549.6 393.46 L575.53 370.92 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M575.53 370.92 L601.49 390.81 L603.61 419.04 L571.04 434.9 L553.34 428.25 L549.6 393.46 L575.53 370.92 Z"
      /><path d="M575.53 370.92 L601.49 390.81 L603.61 419.04 L571.04 434.9 L553.34 428.25 L549.6 393.46 L575.53 370.92 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1044.47 128.92 L1081.42 130.1 L1092.24 149.06 L1080.6801 173.93 L1070.17 178.46 L1035.97 154.78 L1038 136.43 L1044.47 128.92 Z"
      /><path d="M1044.47 128.92 L1081.42 130.1 L1092.24 149.06 L1080.6801 173.93 L1070.17 178.46 L1035.97 154.78 L1038 136.43 L1044.47 128.92 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1044.47 128.92 L1081.42 130.1 L1092.24 149.06 L1080.6801 173.93 L1070.17 178.46 L1035.97 154.78 L1038 136.43 L1044.47 128.92 Z"
      /><path d="M1044.47 128.92 L1081.42 130.1 L1092.24 149.06 L1080.6801 173.93 L1070.17 178.46 L1035.97 154.78 L1038 136.43 L1044.47 128.92 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1044.47 128.92 L1081.42 130.1 L1092.24 149.06 L1080.6801 173.93 L1070.17 178.46 L1035.97 154.78 L1038 136.43 L1044.47 128.92 Z"
      /><path d="M1044.47 128.92 L1081.42 130.1 L1092.24 149.06 L1080.6801 173.93 L1070.17 178.46 L1035.97 154.78 L1038 136.43 L1044.47 128.92 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1044.47 128.92 L1081.42 130.1 L1092.24 149.06 L1080.6801 173.93 L1070.17 178.46 L1035.97 154.78 L1038 136.43 L1044.47 128.92 Z"
      /><path d="M1044.47 128.92 L1081.42 130.1 L1092.24 149.06 L1080.6801 173.93 L1070.17 178.46 L1035.97 154.78 L1038 136.43 L1044.47 128.92 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M872.35 939.1 L914.2 944.68 L915.26 970.5 L878.6 993.78 L872.5 990.99 L860.07 961.8 L872.35 939.1 Z"
      /><path d="M872.35 939.1 L914.2 944.68 L915.26 970.5 L878.6 993.78 L872.5 990.99 L860.07 961.8 L872.35 939.1 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1183.08 194.23 L1167.9 164.4 L1137.1801 168.66 L1127.17 196.34 L1170.8 215.28 L1183.08 194.23 Z"
      /><path d="M1183.08 194.23 L1167.9 164.4 L1137.1801 168.66 L1127.17 196.34 L1170.8 215.28 L1183.08 194.23 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1183.08 194.23 L1167.9 164.4 L1137.1801 168.66 L1127.17 196.34 L1170.8 215.28 L1183.08 194.23 Z"
      /><path d="M1183.08 194.23 L1167.9 164.4 L1137.1801 168.66 L1127.17 196.34 L1170.8 215.28 L1183.08 194.23 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1270.35 783.27 L1230.4 791.58 L1227.92 828.96 L1230.13 831.05 L1274.58 833.23 L1289.9 814.35 L1270.35 783.27 Z"
      /><path d="M1270.35 783.27 L1230.4 791.58 L1227.92 828.96 L1230.13 831.05 L1274.58 833.23 L1289.9 814.35 L1270.35 783.27 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1270.35 783.27 L1230.4 791.58 L1227.92 828.96 L1230.13 831.05 L1274.58 833.23 L1289.9 814.35 L1270.35 783.27 Z"
      /><path d="M1270.35 783.27 L1230.4 791.58 L1227.92 828.96 L1230.13 831.05 L1274.58 833.23 L1289.9 814.35 L1270.35 783.27 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1100.0601 894.58 L1075.4301 927.39 L1091.21 945.14 L1133.1899 934.15 L1133.7 932.8 L1119.51 898.27 L1100.0601 894.58 Z"
      /><path d="M1100.0601 894.58 L1075.4301 927.39 L1091.21 945.14 L1133.1899 934.15 L1133.7 932.8 L1119.51 898.27 L1100.0601 894.58 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1100.0601 894.58 L1075.4301 927.39 L1091.21 945.14 L1133.1899 934.15 L1133.7 932.8 L1119.51 898.27 L1100.0601 894.58 Z"
      /><path d="M1100.0601 894.58 L1075.4301 927.39 L1091.21 945.14 L1133.1899 934.15 L1133.7 932.8 L1119.51 898.27 L1100.0601 894.58 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M815.87 138.01 L795.5 129.14 L771.29 159.63 L782.12 175.02 L820.51 165.31 L815.87 138.01 Z"
      /><path d="M815.87 138.01 L795.5 129.14 L771.29 159.63 L782.12 175.02 L820.51 165.31 L815.87 138.01 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M585.54 695.16 L604.12 726.32 L587.31 746.73 L550.55 738.73 L543.72 724.37 L563.86 696.82 L585.54 695.16 Z"
      /><path d="M585.54 695.16 L604.12 726.32 L587.31 746.73 L550.55 738.73 L543.72 724.37 L563.86 696.82 L585.54 695.16 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M584.23 646.89 L549.13 651.42 L540.59 663.3 L563.86 696.82 L585.54 695.16 L598.66 674.42 L584.23 646.89 Z"
      /><path d="M584.23 646.89 L549.13 651.42 L540.59 663.3 L563.86 696.82 L585.54 695.16 L598.66 674.42 L584.23 646.89 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M584.23 646.89 L549.13 651.42 L540.59 663.3 L563.86 696.82 L585.54 695.16 L598.66 674.42 L584.23 646.89 Z"
      /><path d="M584.23 646.89 L549.13 651.42 L540.59 663.3 L563.86 696.82 L585.54 695.16 L598.66 674.42 L584.23 646.89 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1353.65 708.31 L1365.7 740.73 L1359.77 751.15 L1325.1801 761.94 L1310.14 750.49 L1311.9 720.43 L1344.97 703.61 L1353.65 708.31 Z"
      /><path d="M1353.65 708.31 L1365.7 740.73 L1359.77 751.15 L1325.1801 761.94 L1310.14 750.49 L1311.9 720.43 L1344.97 703.61 L1353.65 708.31 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1353.65 708.31 L1365.7 740.73 L1359.77 751.15 L1325.1801 761.94 L1310.14 750.49 L1311.9 720.43 L1344.97 703.61 L1353.65 708.31 Z"
      /><path d="M1353.65 708.31 L1365.7 740.73 L1359.77 751.15 L1325.1801 761.94 L1310.14 750.49 L1311.9 720.43 L1344.97 703.61 L1353.65 708.31 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1134.52 122.63 L1122.88 147.29 L1137.1801 168.66 L1167.9 164.4 L1177.91 146.08 L1164.64 124.03 L1134.52 122.63 Z"
      /><path d="M1134.52 122.63 L1122.88 147.29 L1137.1801 168.66 L1167.9 164.4 L1177.91 146.08 L1164.64 124.03 L1134.52 122.63 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M582.98 305.27 L590.12 305.37 L612.88 329.98 L575.42 369.03 L551.09 337.73 L582.98 305.27 Z"
      /><path d="M582.98 305.27 L590.12 305.37 L612.88 329.98 L575.42 369.03 L551.09 337.73 L582.98 305.27 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1271.65 191.72 L1253.75 172.39 L1221.03 181.57 L1216.65 188.6 L1230.9 230.56 L1242.95 231.69 L1267.59 215.7 L1271.65 191.72 Z"
      /><path d="M1271.65 191.72 L1253.75 172.39 L1221.03 181.57 L1216.65 188.6 L1230.9 230.56 L1242.95 231.69 L1267.59 215.7 L1271.65 191.72 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1075.4301 927.39 L1061.53 926.05 L1035.45 961.97 L1042.24 976.05 L1072.5601 985.78 L1090.62 969.22 L1091.21 945.14 L1075.4301 927.39 Z"
      /><path d="M1075.4301 927.39 L1061.53 926.05 L1035.45 961.97 L1042.24 976.05 L1072.5601 985.78 L1090.62 969.22 L1091.21 945.14 L1075.4301 927.39 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1075.4301 927.39 L1061.53 926.05 L1035.45 961.97 L1042.24 976.05 L1072.5601 985.78 L1090.62 969.22 L1091.21 945.14 L1075.4301 927.39 Z"
      /><path d="M1075.4301 927.39 L1061.53 926.05 L1035.45 961.97 L1042.24 976.05 L1072.5601 985.78 L1090.62 969.22 L1091.21 945.14 L1075.4301 927.39 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M689.93 254.6 L644.06 234.27 L621.86 262.32 L654.94 298.62 L687.27 278.18 L689.93 254.6 Z"
      /><path d="M689.93 254.6 L644.06 234.27 L621.86 262.32 L654.94 298.62 L687.27 278.18 L689.93 254.6 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M689.93 254.6 L644.06 234.27 L621.86 262.32 L654.94 298.62 L687.27 278.18 L689.93 254.6 Z"
      /><path d="M689.93 254.6 L644.06 234.27 L621.86 262.32 L654.94 298.62 L687.27 278.18 L689.93 254.6 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1213.75 886.6 L1196.05 880.8 L1170.33 899.13 L1169.4 917.75 L1187.84 934.68 L1217.38 920.1 L1213.75 886.6 Z"
      /><path d="M1213.75 886.6 L1196.05 880.8 L1170.33 899.13 L1169.4 917.75 L1187.84 934.68 L1217.38 920.1 L1213.75 886.6 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M621.67 726.2 L644.56 755.74 L640.56 769.98 L617.67 783.67 L592.11 770.57 L587.31 746.73 L604.12 726.32 L621.67 726.2 Z"
      /><path d="M621.67 726.2 L644.56 755.74 L640.56 769.98 L617.67 783.67 L592.11 770.57 L587.31 746.73 L604.12 726.32 L621.67 726.2 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M621.67 726.2 L644.56 755.74 L640.56 769.98 L617.67 783.67 L592.11 770.57 L587.31 746.73 L604.12 726.32 L621.67 726.2 Z"
      /><path d="M621.67 726.2 L644.56 755.74 L640.56 769.98 L617.67 783.67 L592.11 770.57 L587.31 746.73 L604.12 726.32 L621.67 726.2 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M621.67 726.2 L644.56 755.74 L640.56 769.98 L617.67 783.67 L592.11 770.57 L587.31 746.73 L604.12 726.32 L621.67 726.2 Z"
      /><path d="M621.67 726.2 L644.56 755.74 L640.56 769.98 L617.67 783.67 L592.11 770.57 L587.31 746.73 L604.12 726.32 L621.67 726.2 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1230.9 230.56 L1219.04 239.61 L1172.9 230.44 L1170.8 215.28 L1183.08 194.23 L1216.65 188.6 L1230.9 230.56 Z"
      /><path d="M1230.9 230.56 L1219.04 239.61 L1172.9 230.44 L1170.8 215.28 L1183.08 194.23 L1216.65 188.6 L1230.9 230.56 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1230.9 230.56 L1219.04 239.61 L1172.9 230.44 L1170.8 215.28 L1183.08 194.23 L1216.65 188.6 L1230.9 230.56 Z"
      /><path d="M1230.9 230.56 L1219.04 239.61 L1172.9 230.44 L1170.8 215.28 L1183.08 194.23 L1216.65 188.6 L1230.9 230.56 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1230.9 230.56 L1219.04 239.61 L1172.9 230.44 L1170.8 215.28 L1183.08 194.23 L1216.65 188.6 L1230.9 230.56 Z"
      /><path d="M1230.9 230.56 L1219.04 239.61 L1172.9 230.44 L1170.8 215.28 L1183.08 194.23 L1216.65 188.6 L1230.9 230.56 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M706.89 148.93 L729.47 170.58 L726.75 198.67 L707.76 211.4 L673.51 192.33 L674.77 157.64 L689.01 147.67 L706.89 148.93 Z"
      /><path d="M706.89 148.93 L729.47 170.58 L726.75 198.67 L707.76 211.4 L673.51 192.33 L674.77 157.64 L689.01 147.67 L706.89 148.93 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1377.53 629.47 L1338.09 626.6 L1332.53 633.94 L1336.8101 668.87 L1337.3101 669.32 L1387.15 658.52 L1377.53 629.47 Z"
      /><path d="M1377.53 629.47 L1338.09 626.6 L1332.53 633.94 L1336.8101 668.87 L1337.3101 669.32 L1387.15 658.52 L1377.53 629.47 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1377.53 629.47 L1338.09 626.6 L1332.53 633.94 L1336.8101 668.87 L1337.3101 669.32 L1387.15 658.52 L1377.53 629.47 Z"
      /><path d="M1377.53 629.47 L1338.09 626.6 L1332.53 633.94 L1336.8101 668.87 L1337.3101 669.32 L1387.15 658.52 L1377.53 629.47 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1377.53 629.47 L1338.09 626.6 L1332.53 633.94 L1336.8101 668.87 L1337.3101 669.32 L1387.15 658.52 L1377.53 629.47 Z"
      /><path d="M1377.53 629.47 L1338.09 626.6 L1332.53 633.94 L1336.8101 668.87 L1337.3101 669.32 L1387.15 658.52 L1377.53 629.47 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1391.21 661.61 L1387.15 658.52 L1337.3101 669.32 L1344.97 703.61 L1353.65 708.31 L1389.28 691.76 L1391.21 661.61 Z"
      /><path d="M1391.21 661.61 L1387.15 658.52 L1337.3101 669.32 L1344.97 703.61 L1353.65 708.31 L1389.28 691.76 L1391.21 661.61 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M861.92 111.23 L893.5 134.16 L891.65 146.96 L869.9 161.34 L857.65 157.14 L845.53 121.23 L861.92 111.23 Z"
      /><path d="M861.92 111.23 L893.5 134.16 L891.65 146.96 L869.9 161.34 L857.65 157.14 L845.53 121.23 L861.92 111.23 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M861.92 111.23 L893.5 134.16 L891.65 146.96 L869.9 161.34 L857.65 157.14 L845.53 121.23 L861.92 111.23 Z"
      /><path d="M861.92 111.23 L893.5 134.16 L891.65 146.96 L869.9 161.34 L857.65 157.14 L845.53 121.23 L861.92 111.23 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1297.21 266.75 L1264.74 269.07 L1246.76 290.96 L1250.73 314.49 L1269.7 324.31 L1300.3101 306.44 L1300.01 269.75 L1297.21 266.75 Z"
      /><path d="M1297.21 266.75 L1264.74 269.07 L1246.76 290.96 L1250.73 314.49 L1269.7 324.31 L1300.3101 306.44 L1300.01 269.75 L1297.21 266.75 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1297.21 266.75 L1264.74 269.07 L1246.76 290.96 L1250.73 314.49 L1269.7 324.31 L1300.3101 306.44 L1300.01 269.75 L1297.21 266.75 Z"
      /><path d="M1297.21 266.75 L1264.74 269.07 L1246.76 290.96 L1250.73 314.49 L1269.7 324.31 L1300.3101 306.44 L1300.01 269.75 L1297.21 266.75 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1297.21 266.75 L1264.74 269.07 L1246.76 290.96 L1250.73 314.49 L1269.7 324.31 L1300.3101 306.44 L1300.01 269.75 L1297.21 266.75 Z"
      /><path d="M1297.21 266.75 L1264.74 269.07 L1246.76 290.96 L1250.73 314.49 L1269.7 324.31 L1300.3101 306.44 L1300.01 269.75 L1297.21 266.75 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1297.21 266.75 L1264.74 269.07 L1246.76 290.96 L1250.73 314.49 L1269.7 324.31 L1300.3101 306.44 L1300.01 269.75 L1297.21 266.75 Z"
      /><path d="M1297.21 266.75 L1264.74 269.07 L1246.76 290.96 L1250.73 314.49 L1269.7 324.31 L1300.3101 306.44 L1300.01 269.75 L1297.21 266.75 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M989.56 116.82 L971.65 107.1 L950.05 111.25 L937.75 128.48 L943.1 152.5 L959.34 161.09 L985.09 143.44 L990.54 119.73 L989.56 116.82 Z"
      /><path d="M989.56 116.82 L971.65 107.1 L950.05 111.25 L937.75 128.48 L943.1 152.5 L959.34 161.09 L985.09 143.44 L990.54 119.73 L989.56 116.82 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M989.56 116.82 L971.65 107.1 L950.05 111.25 L937.75 128.48 L943.1 152.5 L959.34 161.09 L985.09 143.44 L990.54 119.73 L989.56 116.82 Z"
      /><path d="M989.56 116.82 L971.65 107.1 L950.05 111.25 L937.75 128.48 L943.1 152.5 L959.34 161.09 L985.09 143.44 L990.54 119.73 L989.56 116.82 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M989.56 116.82 L971.65 107.1 L950.05 111.25 L937.75 128.48 L943.1 152.5 L959.34 161.09 L985.09 143.44 L990.54 119.73 L989.56 116.82 Z"
      /><path d="M989.56 116.82 L971.65 107.1 L950.05 111.25 L937.75 128.48 L943.1 152.5 L959.34 161.09 L985.09 143.44 L990.54 119.73 L989.56 116.82 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1404.45 537.68 L1403.91 540.07 L1369.59 557.15 L1352.8101 547.97 L1344.66 515.81 L1380.76 501.69 L1404.45 537.68 Z"
      /><path d="M1404.45 537.68 L1403.91 540.07 L1369.59 557.15 L1352.8101 547.97 L1344.66 515.81 L1380.76 501.69 L1404.45 537.68 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1404.45 537.68 L1403.91 540.07 L1369.59 557.15 L1352.8101 547.97 L1344.66 515.81 L1380.76 501.69 L1404.45 537.68 Z"
      /><path d="M1404.45 537.68 L1403.91 540.07 L1369.59 557.15 L1352.8101 547.97 L1344.66 515.81 L1380.76 501.69 L1404.45 537.68 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1404.45 537.68 L1403.91 540.07 L1369.59 557.15 L1352.8101 547.97 L1344.66 515.81 L1380.76 501.69 L1404.45 537.68 Z"
      /><path d="M1404.45 537.68 L1403.91 540.07 L1369.59 557.15 L1352.8101 547.97 L1344.66 515.81 L1380.76 501.69 L1404.45 537.68 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1350.8 270.86 L1300.01 269.75 L1300.3101 306.44 L1330.4301 324.89 L1342.34 320.92 L1350.8 270.86 Z"
      /><path d="M1350.8 270.86 L1300.01 269.75 L1300.3101 306.44 L1330.4301 324.89 L1342.34 320.92 L1350.8 270.86 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M971 913.61 L955.65 935.97 L973.36 970.28 L981.79 972.02 L1011.13 953.43 L1003.63 913.93 L971 913.61 Z"
      /><path d="M971 913.61 L955.65 935.97 L973.36 970.28 L981.79 972.02 L1011.13 953.43 L1003.63 913.93 L971 913.61 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M971 913.61 L955.65 935.97 L973.36 970.28 L981.79 972.02 L1011.13 953.43 L1003.63 913.93 L971 913.61 Z"
      /><path d="M971 913.61 L955.65 935.97 L973.36 970.28 L981.79 972.02 L1011.13 953.43 L1003.63 913.93 L971 913.61 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M971 913.61 L955.65 935.97 L973.36 970.28 L981.79 972.02 L1011.13 953.43 L1003.63 913.93 L971 913.61 Z"
      /><path d="M971 913.61 L955.65 935.97 L973.36 970.28 L981.79 972.02 L1011.13 953.43 L1003.63 913.93 L971 913.61 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M708.1 839.98 L713.54 865.6 L674.67 881.7 L653.25 862.29 L660.31 827.04 L666.53 822.38 L708.1 839.98 Z"
      /><path d="M708.1 839.98 L713.54 865.6 L674.67 881.7 L653.25 862.29 L660.31 827.04 L666.53 822.38 L708.1 839.98 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M708.1 839.98 L713.54 865.6 L674.67 881.7 L653.25 862.29 L660.31 827.04 L666.53 822.38 L708.1 839.98 Z"
      /><path d="M708.1 839.98 L713.54 865.6 L674.67 881.7 L653.25 862.29 L660.31 827.04 L666.53 822.38 L708.1 839.98 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1370.6801 333.49 L1342.34 320.92 L1330.4301 324.89 L1314.8 360.56 L1321.41 375.04 L1367.0601 382.52 L1370.6801 333.49 Z"
      /><path d="M1370.6801 333.49 L1342.34 320.92 L1330.4301 324.89 L1314.8 360.56 L1321.41 375.04 L1367.0601 382.52 L1370.6801 333.49 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1370.6801 333.49 L1342.34 320.92 L1330.4301 324.89 L1314.8 360.56 L1321.41 375.04 L1367.0601 382.52 L1370.6801 333.49 Z"
      /><path d="M1370.6801 333.49 L1342.34 320.92 L1330.4301 324.89 L1314.8 360.56 L1321.41 375.04 L1367.0601 382.52 L1370.6801 333.49 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M845.53 121.23 L857.65 157.14 L828.67 171.16 L820.51 165.31 L815.87 138.01 L841.19 120.69 L845.53 121.23 Z"
      /><path d="M845.53 121.23 L857.65 157.14 L828.67 171.16 L820.51 165.31 L815.87 138.01 L841.19 120.69 L845.53 121.23 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M845.53 121.23 L857.65 157.14 L828.67 171.16 L820.51 165.31 L815.87 138.01 L841.19 120.69 L845.53 121.23 Z"
      /><path d="M845.53 121.23 L857.65 157.14 L828.67 171.16 L820.51 165.31 L815.87 138.01 L841.19 120.69 L845.53 121.23 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M545.94 491.11 L523.99 523.57 L546.29 553.73 L549.36 553.89 L576.22 530.26 L558.18 491.95 L545.94 491.11 Z"
      /><path d="M545.94 491.11 L523.99 523.57 L546.29 553.73 L549.36 553.89 L576.22 530.26 L558.18 491.95 L545.94 491.11 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M545.94 491.11 L523.99 523.57 L546.29 553.73 L549.36 553.89 L576.22 530.26 L558.18 491.95 L545.94 491.11 Z"
      /><path d="M545.94 491.11 L523.99 523.57 L546.29 553.73 L549.36 553.89 L576.22 530.26 L558.18 491.95 L545.94 491.11 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M543.75 336.54 L551.09 337.73 L575.42 369.03 L575.53 370.92 L549.6 393.46 L516.64 381.26 L520.45 351.88 L543.75 336.54 Z"
      /><path d="M543.75 336.54 L551.09 337.73 L575.42 369.03 L575.53 370.92 L549.6 393.46 L516.64 381.26 L520.45 351.88 L543.75 336.54 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1106.1 96.92 L1125.02 103.95 L1134.52 122.63 L1122.88 147.29 L1092.24 149.06 L1081.42 130.1 L1091.0601 103.39 L1106.1 96.92 Z"
      /><path d="M1106.1 96.92 L1125.02 103.95 L1134.52 122.63 L1122.88 147.29 L1092.24 149.06 L1081.42 130.1 L1091.0601 103.39 L1106.1 96.92 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M707.76 211.4 L704.5 242.05 L689.93 254.6 L644.06 234.27 L642.48 212.11 L673.51 192.33 L707.76 211.4 Z"
      /><path d="M707.76 211.4 L704.5 242.05 L689.93 254.6 L644.06 234.27 L642.48 212.11 L673.51 192.33 L707.76 211.4 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M707.76 211.4 L704.5 242.05 L689.93 254.6 L644.06 234.27 L642.48 212.11 L673.51 192.33 L707.76 211.4 Z"
      /><path d="M707.76 211.4 L704.5 242.05 L689.93 254.6 L644.06 234.27 L642.48 212.11 L673.51 192.33 L707.76 211.4 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1310.14 750.49 L1325.1801 761.94 L1327 792.95 L1305.04 814.21 L1289.9 814.35 L1270.35 783.27 L1277.4301 760.51 L1310.14 750.49 Z"
      /><path d="M1310.14 750.49 L1325.1801 761.94 L1327 792.95 L1305.04 814.21 L1289.9 814.35 L1270.35 783.27 L1277.4301 760.51 L1310.14 750.49 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1310.14 750.49 L1325.1801 761.94 L1327 792.95 L1305.04 814.21 L1289.9 814.35 L1270.35 783.27 L1277.4301 760.51 L1310.14 750.49 Z"
      /><path d="M1310.14 750.49 L1325.1801 761.94 L1327 792.95 L1305.04 814.21 L1289.9 814.35 L1270.35 783.27 L1277.4301 760.51 L1310.14 750.49 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M760.31 156.27 L771.29 159.63 L782.12 175.02 L781.08 195.16 L758.09 212.02 L726.75 198.67 L729.47 170.58 L760.31 156.27 Z"
      /><path d="M760.31 156.27 L771.29 159.63 L782.12 175.02 L781.08 195.16 L758.09 212.02 L726.75 198.67 L729.47 170.58 L760.31 156.27 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M760.31 156.27 L771.29 159.63 L782.12 175.02 L781.08 195.16 L758.09 212.02 L726.75 198.67 L729.47 170.58 L760.31 156.27 Z"
      /><path d="M760.31 156.27 L771.29 159.63 L782.12 175.02 L781.08 195.16 L758.09 212.02 L726.75 198.67 L729.47 170.58 L760.31 156.27 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M760.31 156.27 L771.29 159.63 L782.12 175.02 L781.08 195.16 L758.09 212.02 L726.75 198.67 L729.47 170.58 L760.31 156.27 Z"
      /><path d="M760.31 156.27 L771.29 159.63 L782.12 175.02 L781.08 195.16 L758.09 212.02 L726.75 198.67 L729.47 170.58 L760.31 156.27 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1299.6 236.39 L1297.21 266.75 L1264.74 269.07 L1242.95 231.69 L1267.59 215.7 L1299.6 236.39 Z"
      /><path d="M1299.6 236.39 L1297.21 266.75 L1264.74 269.07 L1242.95 231.69 L1267.59 215.7 L1299.6 236.39 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M937.75 128.48 L907.38 121.6 L893.5 134.16 L891.65 146.96 L916.46 167.32 L943.1 152.5 L937.75 128.48 Z"
      /><path d="M937.75 128.48 L907.38 121.6 L893.5 134.16 L891.65 146.96 L916.46 167.32 L943.1 152.5 L937.75 128.48 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M937.75 128.48 L907.38 121.6 L893.5 134.16 L891.65 146.96 L916.46 167.32 L943.1 152.5 L937.75 128.48 Z"
      /><path d="M937.75 128.48 L907.38 121.6 L893.5 134.16 L891.65 146.96 L916.46 167.32 L943.1 152.5 L937.75 128.48 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1370.8101 585.77 L1391.3 602.91 L1377.53 629.47 L1338.09 626.6 L1336.17 598.08 L1370.8101 585.77 Z"
      /><path d="M1370.8101 585.77 L1391.3 602.91 L1377.53 629.47 L1338.09 626.6 L1336.17 598.08 L1370.8101 585.77 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1370.8101 585.77 L1391.3 602.91 L1377.53 629.47 L1338.09 626.6 L1336.17 598.08 L1370.8101 585.77 Z"
      /><path d="M1370.8101 585.77 L1391.3 602.91 L1377.53 629.47 L1338.09 626.6 L1336.17 598.08 L1370.8101 585.77 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M776.43 886.29 L810.8 890.77 L820.83 918.6 L812.13 935.41 L773 939.25 L761.68 907.08 L776.43 886.29 Z"
      /><path d="M776.43 886.29 L810.8 890.77 L820.83 918.6 L812.13 935.41 L773 939.25 L761.68 907.08 L776.43 886.29 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M776.43 886.29 L810.8 890.77 L820.83 918.6 L812.13 935.41 L773 939.25 L761.68 907.08 L776.43 886.29 Z"
      /><path d="M776.43 886.29 L810.8 890.77 L820.83 918.6 L812.13 935.41 L773 939.25 L761.68 907.08 L776.43 886.29 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1230.13 831.05 L1227.92 828.96 L1189.52 834.64 L1183.55 849 L1196.05 880.8 L1213.75 886.6 L1233.39 874.91 L1230.13 831.05 Z"
      /><path d="M1230.13 831.05 L1227.92 828.96 L1189.52 834.64 L1183.55 849 L1196.05 880.8 L1213.75 886.6 L1233.39 874.91 L1230.13 831.05 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1230.13 831.05 L1227.92 828.96 L1189.52 834.64 L1183.55 849 L1196.05 880.8 L1213.75 886.6 L1233.39 874.91 L1230.13 831.05 Z"
      /><path d="M1230.13 831.05 L1227.92 828.96 L1189.52 834.64 L1183.55 849 L1196.05 880.8 L1213.75 886.6 L1233.39 874.91 L1230.13 831.05 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1230.13 831.05 L1227.92 828.96 L1189.52 834.64 L1183.55 849 L1196.05 880.8 L1213.75 886.6 L1233.39 874.91 L1230.13 831.05 Z"
      /><path d="M1230.13 831.05 L1227.92 828.96 L1189.52 834.64 L1183.55 849 L1196.05 880.8 L1213.75 886.6 L1233.39 874.91 L1230.13 831.05 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M654.94 298.62 L621.86 262.32 L615.46 263.35 L590.12 305.37 L612.88 329.98 L617.62 331.02 L652.81 310.23 L654.94 298.62 Z"
      /><path d="M654.94 298.62 L621.86 262.32 L615.46 263.35 L590.12 305.37 L612.88 329.98 L617.62 331.02 L652.81 310.23 L654.94 298.62 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M654.94 298.62 L621.86 262.32 L615.46 263.35 L590.12 305.37 L612.88 329.98 L617.62 331.02 L652.81 310.23 L654.94 298.62 Z"
      /><path d="M654.94 298.62 L621.86 262.32 L615.46 263.35 L590.12 305.37 L612.88 329.98 L617.62 331.02 L652.81 310.23 L654.94 298.62 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M654.94 298.62 L621.86 262.32 L615.46 263.35 L590.12 305.37 L612.88 329.98 L617.62 331.02 L652.81 310.23 L654.94 298.62 Z"
      /><path d="M654.94 298.62 L621.86 262.32 L615.46 263.35 L590.12 305.37 L612.88 329.98 L617.62 331.02 L652.81 310.23 L654.94 298.62 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1418.89 564.96 L1403.91 540.07 L1369.59 557.15 L1370.8101 585.77 L1391.3 602.91 L1398.9399 601.52 L1418.89 564.96 Z"
      /><path d="M1418.89 564.96 L1403.91 540.07 L1369.59 557.15 L1370.8101 585.77 L1391.3 602.91 L1398.9399 601.52 L1418.89 564.96 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M1035.45 961.97 L1011.13 953.43 L981.79 972.02 L1001.66 1012.65 L1020.45 1013.34 L1042.24 976.05 L1035.45 961.97 Z"
      /><path d="M1035.45 961.97 L1011.13 953.43 L981.79 972.02 L1001.66 1012.65 L1020.45 1013.34 L1042.24 976.05 L1035.45 961.97 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M571.96 599.49 L540.07 613.4 L549.13 651.42 L584.23 646.89 L593.45 627.44 L571.96 599.49 Z"
      /><path d="M571.96 599.49 L540.07 613.4 L549.13 651.42 L584.23 646.89 L593.45 627.44 L571.96 599.49 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M571.96 599.49 L540.07 613.4 L549.13 651.42 L584.23 646.89 L593.45 627.44 L571.96 599.49 Z"
      /><path d="M571.96 599.49 L540.07 613.4 L549.13 651.42 L584.23 646.89 L593.45 627.44 L571.96 599.49 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M776.43 886.29 L766.24 855.73 L714.68 866.34 L728.43 904.21 L761.68 907.08 L776.43 886.29 Z"
      /><path d="M776.43 886.29 L766.24 855.73 L714.68 866.34 L728.43 904.21 L761.68 907.08 L776.43 886.29 Z" style="fill:rgb(47,177,0); stroke:none;"
      /><path style="fill:none;" d="M776.43 886.29 L766.24 855.73 L714.68 866.34 L728.43 904.21 L761.68 907.08 L776.43 886.29 Z"
      /><path d="M776.43 886.29 L766.24 855.73 L714.68 866.34 L728.43 904.21 L761.68 907.08 L776.43 886.29 Z" style="fill:rgb(47,177,0); stroke:none;"
    /></g
  ></g
></svg
>
